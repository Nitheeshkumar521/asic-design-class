module RV_CPU (clk,
    reset,
    out);
 input clk;
 input reset;
 output [9:0] out;

 wire \CPU_Dmem_value_a5[0][0] ;
 wire \CPU_Dmem_value_a5[0][10] ;
 wire \CPU_Dmem_value_a5[0][11] ;
 wire \CPU_Dmem_value_a5[0][12] ;
 wire \CPU_Dmem_value_a5[0][13] ;
 wire \CPU_Dmem_value_a5[0][14] ;
 wire \CPU_Dmem_value_a5[0][15] ;
 wire \CPU_Dmem_value_a5[0][16] ;
 wire \CPU_Dmem_value_a5[0][17] ;
 wire \CPU_Dmem_value_a5[0][18] ;
 wire \CPU_Dmem_value_a5[0][19] ;
 wire \CPU_Dmem_value_a5[0][1] ;
 wire \CPU_Dmem_value_a5[0][20] ;
 wire \CPU_Dmem_value_a5[0][21] ;
 wire \CPU_Dmem_value_a5[0][22] ;
 wire \CPU_Dmem_value_a5[0][23] ;
 wire \CPU_Dmem_value_a5[0][24] ;
 wire \CPU_Dmem_value_a5[0][25] ;
 wire \CPU_Dmem_value_a5[0][26] ;
 wire \CPU_Dmem_value_a5[0][27] ;
 wire \CPU_Dmem_value_a5[0][28] ;
 wire \CPU_Dmem_value_a5[0][29] ;
 wire \CPU_Dmem_value_a5[0][2] ;
 wire \CPU_Dmem_value_a5[0][30] ;
 wire \CPU_Dmem_value_a5[0][31] ;
 wire \CPU_Dmem_value_a5[0][3] ;
 wire \CPU_Dmem_value_a5[0][4] ;
 wire \CPU_Dmem_value_a5[0][5] ;
 wire \CPU_Dmem_value_a5[0][6] ;
 wire \CPU_Dmem_value_a5[0][7] ;
 wire \CPU_Dmem_value_a5[0][8] ;
 wire \CPU_Dmem_value_a5[0][9] ;
 wire \CPU_Dmem_value_a5[10][0] ;
 wire \CPU_Dmem_value_a5[10][10] ;
 wire \CPU_Dmem_value_a5[10][11] ;
 wire \CPU_Dmem_value_a5[10][12] ;
 wire \CPU_Dmem_value_a5[10][13] ;
 wire \CPU_Dmem_value_a5[10][14] ;
 wire \CPU_Dmem_value_a5[10][15] ;
 wire \CPU_Dmem_value_a5[10][16] ;
 wire \CPU_Dmem_value_a5[10][17] ;
 wire \CPU_Dmem_value_a5[10][18] ;
 wire \CPU_Dmem_value_a5[10][19] ;
 wire \CPU_Dmem_value_a5[10][1] ;
 wire \CPU_Dmem_value_a5[10][20] ;
 wire \CPU_Dmem_value_a5[10][21] ;
 wire \CPU_Dmem_value_a5[10][22] ;
 wire \CPU_Dmem_value_a5[10][23] ;
 wire \CPU_Dmem_value_a5[10][24] ;
 wire \CPU_Dmem_value_a5[10][25] ;
 wire \CPU_Dmem_value_a5[10][26] ;
 wire \CPU_Dmem_value_a5[10][27] ;
 wire \CPU_Dmem_value_a5[10][28] ;
 wire \CPU_Dmem_value_a5[10][29] ;
 wire \CPU_Dmem_value_a5[10][2] ;
 wire \CPU_Dmem_value_a5[10][30] ;
 wire \CPU_Dmem_value_a5[10][31] ;
 wire \CPU_Dmem_value_a5[10][3] ;
 wire \CPU_Dmem_value_a5[10][4] ;
 wire \CPU_Dmem_value_a5[10][5] ;
 wire \CPU_Dmem_value_a5[10][6] ;
 wire \CPU_Dmem_value_a5[10][7] ;
 wire \CPU_Dmem_value_a5[10][8] ;
 wire \CPU_Dmem_value_a5[10][9] ;
 wire \CPU_Dmem_value_a5[11][0] ;
 wire \CPU_Dmem_value_a5[11][10] ;
 wire \CPU_Dmem_value_a5[11][11] ;
 wire \CPU_Dmem_value_a5[11][12] ;
 wire \CPU_Dmem_value_a5[11][13] ;
 wire \CPU_Dmem_value_a5[11][14] ;
 wire \CPU_Dmem_value_a5[11][15] ;
 wire \CPU_Dmem_value_a5[11][16] ;
 wire \CPU_Dmem_value_a5[11][17] ;
 wire \CPU_Dmem_value_a5[11][18] ;
 wire \CPU_Dmem_value_a5[11][19] ;
 wire \CPU_Dmem_value_a5[11][1] ;
 wire \CPU_Dmem_value_a5[11][20] ;
 wire \CPU_Dmem_value_a5[11][21] ;
 wire \CPU_Dmem_value_a5[11][22] ;
 wire \CPU_Dmem_value_a5[11][23] ;
 wire \CPU_Dmem_value_a5[11][24] ;
 wire \CPU_Dmem_value_a5[11][25] ;
 wire \CPU_Dmem_value_a5[11][26] ;
 wire \CPU_Dmem_value_a5[11][27] ;
 wire \CPU_Dmem_value_a5[11][28] ;
 wire \CPU_Dmem_value_a5[11][29] ;
 wire \CPU_Dmem_value_a5[11][2] ;
 wire \CPU_Dmem_value_a5[11][30] ;
 wire \CPU_Dmem_value_a5[11][31] ;
 wire \CPU_Dmem_value_a5[11][3] ;
 wire \CPU_Dmem_value_a5[11][4] ;
 wire \CPU_Dmem_value_a5[11][5] ;
 wire \CPU_Dmem_value_a5[11][6] ;
 wire \CPU_Dmem_value_a5[11][7] ;
 wire \CPU_Dmem_value_a5[11][8] ;
 wire \CPU_Dmem_value_a5[11][9] ;
 wire \CPU_Dmem_value_a5[12][0] ;
 wire \CPU_Dmem_value_a5[12][10] ;
 wire \CPU_Dmem_value_a5[12][11] ;
 wire \CPU_Dmem_value_a5[12][12] ;
 wire \CPU_Dmem_value_a5[12][13] ;
 wire \CPU_Dmem_value_a5[12][14] ;
 wire \CPU_Dmem_value_a5[12][15] ;
 wire \CPU_Dmem_value_a5[12][16] ;
 wire \CPU_Dmem_value_a5[12][17] ;
 wire \CPU_Dmem_value_a5[12][18] ;
 wire \CPU_Dmem_value_a5[12][19] ;
 wire \CPU_Dmem_value_a5[12][1] ;
 wire \CPU_Dmem_value_a5[12][20] ;
 wire \CPU_Dmem_value_a5[12][21] ;
 wire \CPU_Dmem_value_a5[12][22] ;
 wire \CPU_Dmem_value_a5[12][23] ;
 wire \CPU_Dmem_value_a5[12][24] ;
 wire \CPU_Dmem_value_a5[12][25] ;
 wire \CPU_Dmem_value_a5[12][26] ;
 wire \CPU_Dmem_value_a5[12][27] ;
 wire \CPU_Dmem_value_a5[12][28] ;
 wire \CPU_Dmem_value_a5[12][29] ;
 wire \CPU_Dmem_value_a5[12][2] ;
 wire \CPU_Dmem_value_a5[12][30] ;
 wire \CPU_Dmem_value_a5[12][31] ;
 wire \CPU_Dmem_value_a5[12][3] ;
 wire \CPU_Dmem_value_a5[12][4] ;
 wire \CPU_Dmem_value_a5[12][5] ;
 wire \CPU_Dmem_value_a5[12][6] ;
 wire \CPU_Dmem_value_a5[12][7] ;
 wire \CPU_Dmem_value_a5[12][8] ;
 wire \CPU_Dmem_value_a5[12][9] ;
 wire \CPU_Dmem_value_a5[13][0] ;
 wire \CPU_Dmem_value_a5[13][10] ;
 wire \CPU_Dmem_value_a5[13][11] ;
 wire \CPU_Dmem_value_a5[13][12] ;
 wire \CPU_Dmem_value_a5[13][13] ;
 wire \CPU_Dmem_value_a5[13][14] ;
 wire \CPU_Dmem_value_a5[13][15] ;
 wire \CPU_Dmem_value_a5[13][16] ;
 wire \CPU_Dmem_value_a5[13][17] ;
 wire \CPU_Dmem_value_a5[13][18] ;
 wire \CPU_Dmem_value_a5[13][19] ;
 wire \CPU_Dmem_value_a5[13][1] ;
 wire \CPU_Dmem_value_a5[13][20] ;
 wire \CPU_Dmem_value_a5[13][21] ;
 wire \CPU_Dmem_value_a5[13][22] ;
 wire \CPU_Dmem_value_a5[13][23] ;
 wire \CPU_Dmem_value_a5[13][24] ;
 wire \CPU_Dmem_value_a5[13][25] ;
 wire \CPU_Dmem_value_a5[13][26] ;
 wire \CPU_Dmem_value_a5[13][27] ;
 wire \CPU_Dmem_value_a5[13][28] ;
 wire \CPU_Dmem_value_a5[13][29] ;
 wire \CPU_Dmem_value_a5[13][2] ;
 wire \CPU_Dmem_value_a5[13][30] ;
 wire \CPU_Dmem_value_a5[13][31] ;
 wire \CPU_Dmem_value_a5[13][3] ;
 wire \CPU_Dmem_value_a5[13][4] ;
 wire \CPU_Dmem_value_a5[13][5] ;
 wire \CPU_Dmem_value_a5[13][6] ;
 wire \CPU_Dmem_value_a5[13][7] ;
 wire \CPU_Dmem_value_a5[13][8] ;
 wire \CPU_Dmem_value_a5[13][9] ;
 wire \CPU_Dmem_value_a5[14][0] ;
 wire \CPU_Dmem_value_a5[14][10] ;
 wire \CPU_Dmem_value_a5[14][11] ;
 wire \CPU_Dmem_value_a5[14][12] ;
 wire \CPU_Dmem_value_a5[14][13] ;
 wire \CPU_Dmem_value_a5[14][14] ;
 wire \CPU_Dmem_value_a5[14][15] ;
 wire \CPU_Dmem_value_a5[14][16] ;
 wire \CPU_Dmem_value_a5[14][17] ;
 wire \CPU_Dmem_value_a5[14][18] ;
 wire \CPU_Dmem_value_a5[14][19] ;
 wire \CPU_Dmem_value_a5[14][1] ;
 wire \CPU_Dmem_value_a5[14][20] ;
 wire \CPU_Dmem_value_a5[14][21] ;
 wire \CPU_Dmem_value_a5[14][22] ;
 wire \CPU_Dmem_value_a5[14][23] ;
 wire \CPU_Dmem_value_a5[14][24] ;
 wire \CPU_Dmem_value_a5[14][25] ;
 wire \CPU_Dmem_value_a5[14][26] ;
 wire \CPU_Dmem_value_a5[14][27] ;
 wire \CPU_Dmem_value_a5[14][28] ;
 wire \CPU_Dmem_value_a5[14][29] ;
 wire \CPU_Dmem_value_a5[14][2] ;
 wire \CPU_Dmem_value_a5[14][30] ;
 wire \CPU_Dmem_value_a5[14][31] ;
 wire \CPU_Dmem_value_a5[14][3] ;
 wire \CPU_Dmem_value_a5[14][4] ;
 wire \CPU_Dmem_value_a5[14][5] ;
 wire \CPU_Dmem_value_a5[14][6] ;
 wire \CPU_Dmem_value_a5[14][7] ;
 wire \CPU_Dmem_value_a5[14][8] ;
 wire \CPU_Dmem_value_a5[14][9] ;
 wire \CPU_Dmem_value_a5[15][0] ;
 wire \CPU_Dmem_value_a5[15][10] ;
 wire \CPU_Dmem_value_a5[15][11] ;
 wire \CPU_Dmem_value_a5[15][12] ;
 wire \CPU_Dmem_value_a5[15][13] ;
 wire \CPU_Dmem_value_a5[15][14] ;
 wire \CPU_Dmem_value_a5[15][15] ;
 wire \CPU_Dmem_value_a5[15][16] ;
 wire \CPU_Dmem_value_a5[15][17] ;
 wire \CPU_Dmem_value_a5[15][18] ;
 wire \CPU_Dmem_value_a5[15][19] ;
 wire \CPU_Dmem_value_a5[15][1] ;
 wire \CPU_Dmem_value_a5[15][20] ;
 wire \CPU_Dmem_value_a5[15][21] ;
 wire \CPU_Dmem_value_a5[15][22] ;
 wire \CPU_Dmem_value_a5[15][23] ;
 wire \CPU_Dmem_value_a5[15][24] ;
 wire \CPU_Dmem_value_a5[15][25] ;
 wire \CPU_Dmem_value_a5[15][26] ;
 wire \CPU_Dmem_value_a5[15][27] ;
 wire \CPU_Dmem_value_a5[15][28] ;
 wire \CPU_Dmem_value_a5[15][29] ;
 wire \CPU_Dmem_value_a5[15][2] ;
 wire \CPU_Dmem_value_a5[15][30] ;
 wire \CPU_Dmem_value_a5[15][31] ;
 wire \CPU_Dmem_value_a5[15][3] ;
 wire \CPU_Dmem_value_a5[15][4] ;
 wire \CPU_Dmem_value_a5[15][5] ;
 wire \CPU_Dmem_value_a5[15][6] ;
 wire \CPU_Dmem_value_a5[15][7] ;
 wire \CPU_Dmem_value_a5[15][8] ;
 wire \CPU_Dmem_value_a5[15][9] ;
 wire \CPU_Dmem_value_a5[1][0] ;
 wire \CPU_Dmem_value_a5[1][10] ;
 wire \CPU_Dmem_value_a5[1][11] ;
 wire \CPU_Dmem_value_a5[1][12] ;
 wire \CPU_Dmem_value_a5[1][13] ;
 wire \CPU_Dmem_value_a5[1][14] ;
 wire \CPU_Dmem_value_a5[1][15] ;
 wire \CPU_Dmem_value_a5[1][16] ;
 wire \CPU_Dmem_value_a5[1][17] ;
 wire \CPU_Dmem_value_a5[1][18] ;
 wire \CPU_Dmem_value_a5[1][19] ;
 wire \CPU_Dmem_value_a5[1][1] ;
 wire \CPU_Dmem_value_a5[1][20] ;
 wire \CPU_Dmem_value_a5[1][21] ;
 wire \CPU_Dmem_value_a5[1][22] ;
 wire \CPU_Dmem_value_a5[1][23] ;
 wire \CPU_Dmem_value_a5[1][24] ;
 wire \CPU_Dmem_value_a5[1][25] ;
 wire \CPU_Dmem_value_a5[1][26] ;
 wire \CPU_Dmem_value_a5[1][27] ;
 wire \CPU_Dmem_value_a5[1][28] ;
 wire \CPU_Dmem_value_a5[1][29] ;
 wire \CPU_Dmem_value_a5[1][2] ;
 wire \CPU_Dmem_value_a5[1][30] ;
 wire \CPU_Dmem_value_a5[1][31] ;
 wire \CPU_Dmem_value_a5[1][3] ;
 wire \CPU_Dmem_value_a5[1][4] ;
 wire \CPU_Dmem_value_a5[1][5] ;
 wire \CPU_Dmem_value_a5[1][6] ;
 wire \CPU_Dmem_value_a5[1][7] ;
 wire \CPU_Dmem_value_a5[1][8] ;
 wire \CPU_Dmem_value_a5[1][9] ;
 wire \CPU_Dmem_value_a5[2][0] ;
 wire \CPU_Dmem_value_a5[2][10] ;
 wire \CPU_Dmem_value_a5[2][11] ;
 wire \CPU_Dmem_value_a5[2][12] ;
 wire \CPU_Dmem_value_a5[2][13] ;
 wire \CPU_Dmem_value_a5[2][14] ;
 wire \CPU_Dmem_value_a5[2][15] ;
 wire \CPU_Dmem_value_a5[2][16] ;
 wire \CPU_Dmem_value_a5[2][17] ;
 wire \CPU_Dmem_value_a5[2][18] ;
 wire \CPU_Dmem_value_a5[2][19] ;
 wire \CPU_Dmem_value_a5[2][1] ;
 wire \CPU_Dmem_value_a5[2][20] ;
 wire \CPU_Dmem_value_a5[2][21] ;
 wire \CPU_Dmem_value_a5[2][22] ;
 wire \CPU_Dmem_value_a5[2][23] ;
 wire \CPU_Dmem_value_a5[2][24] ;
 wire \CPU_Dmem_value_a5[2][25] ;
 wire \CPU_Dmem_value_a5[2][26] ;
 wire \CPU_Dmem_value_a5[2][27] ;
 wire \CPU_Dmem_value_a5[2][28] ;
 wire \CPU_Dmem_value_a5[2][29] ;
 wire \CPU_Dmem_value_a5[2][2] ;
 wire \CPU_Dmem_value_a5[2][30] ;
 wire \CPU_Dmem_value_a5[2][31] ;
 wire \CPU_Dmem_value_a5[2][3] ;
 wire \CPU_Dmem_value_a5[2][4] ;
 wire \CPU_Dmem_value_a5[2][5] ;
 wire \CPU_Dmem_value_a5[2][6] ;
 wire \CPU_Dmem_value_a5[2][7] ;
 wire \CPU_Dmem_value_a5[2][8] ;
 wire \CPU_Dmem_value_a5[2][9] ;
 wire \CPU_Dmem_value_a5[3][0] ;
 wire \CPU_Dmem_value_a5[3][10] ;
 wire \CPU_Dmem_value_a5[3][11] ;
 wire \CPU_Dmem_value_a5[3][12] ;
 wire \CPU_Dmem_value_a5[3][13] ;
 wire \CPU_Dmem_value_a5[3][14] ;
 wire \CPU_Dmem_value_a5[3][15] ;
 wire \CPU_Dmem_value_a5[3][16] ;
 wire \CPU_Dmem_value_a5[3][17] ;
 wire \CPU_Dmem_value_a5[3][18] ;
 wire \CPU_Dmem_value_a5[3][19] ;
 wire \CPU_Dmem_value_a5[3][1] ;
 wire \CPU_Dmem_value_a5[3][20] ;
 wire \CPU_Dmem_value_a5[3][21] ;
 wire \CPU_Dmem_value_a5[3][22] ;
 wire \CPU_Dmem_value_a5[3][23] ;
 wire \CPU_Dmem_value_a5[3][24] ;
 wire \CPU_Dmem_value_a5[3][25] ;
 wire \CPU_Dmem_value_a5[3][26] ;
 wire \CPU_Dmem_value_a5[3][27] ;
 wire \CPU_Dmem_value_a5[3][28] ;
 wire \CPU_Dmem_value_a5[3][29] ;
 wire \CPU_Dmem_value_a5[3][2] ;
 wire \CPU_Dmem_value_a5[3][30] ;
 wire \CPU_Dmem_value_a5[3][31] ;
 wire \CPU_Dmem_value_a5[3][3] ;
 wire \CPU_Dmem_value_a5[3][4] ;
 wire \CPU_Dmem_value_a5[3][5] ;
 wire \CPU_Dmem_value_a5[3][6] ;
 wire \CPU_Dmem_value_a5[3][7] ;
 wire \CPU_Dmem_value_a5[3][8] ;
 wire \CPU_Dmem_value_a5[3][9] ;
 wire \CPU_Dmem_value_a5[4][0] ;
 wire \CPU_Dmem_value_a5[4][10] ;
 wire \CPU_Dmem_value_a5[4][11] ;
 wire \CPU_Dmem_value_a5[4][12] ;
 wire \CPU_Dmem_value_a5[4][13] ;
 wire \CPU_Dmem_value_a5[4][14] ;
 wire \CPU_Dmem_value_a5[4][15] ;
 wire \CPU_Dmem_value_a5[4][16] ;
 wire \CPU_Dmem_value_a5[4][17] ;
 wire \CPU_Dmem_value_a5[4][18] ;
 wire \CPU_Dmem_value_a5[4][19] ;
 wire \CPU_Dmem_value_a5[4][1] ;
 wire \CPU_Dmem_value_a5[4][20] ;
 wire \CPU_Dmem_value_a5[4][21] ;
 wire \CPU_Dmem_value_a5[4][22] ;
 wire \CPU_Dmem_value_a5[4][23] ;
 wire \CPU_Dmem_value_a5[4][24] ;
 wire \CPU_Dmem_value_a5[4][25] ;
 wire \CPU_Dmem_value_a5[4][26] ;
 wire \CPU_Dmem_value_a5[4][27] ;
 wire \CPU_Dmem_value_a5[4][28] ;
 wire \CPU_Dmem_value_a5[4][29] ;
 wire \CPU_Dmem_value_a5[4][2] ;
 wire \CPU_Dmem_value_a5[4][30] ;
 wire \CPU_Dmem_value_a5[4][31] ;
 wire \CPU_Dmem_value_a5[4][3] ;
 wire \CPU_Dmem_value_a5[4][4] ;
 wire \CPU_Dmem_value_a5[4][5] ;
 wire \CPU_Dmem_value_a5[4][6] ;
 wire \CPU_Dmem_value_a5[4][7] ;
 wire \CPU_Dmem_value_a5[4][8] ;
 wire \CPU_Dmem_value_a5[4][9] ;
 wire \CPU_Dmem_value_a5[5][0] ;
 wire \CPU_Dmem_value_a5[5][10] ;
 wire \CPU_Dmem_value_a5[5][11] ;
 wire \CPU_Dmem_value_a5[5][12] ;
 wire \CPU_Dmem_value_a5[5][13] ;
 wire \CPU_Dmem_value_a5[5][14] ;
 wire \CPU_Dmem_value_a5[5][15] ;
 wire \CPU_Dmem_value_a5[5][16] ;
 wire \CPU_Dmem_value_a5[5][17] ;
 wire \CPU_Dmem_value_a5[5][18] ;
 wire \CPU_Dmem_value_a5[5][19] ;
 wire \CPU_Dmem_value_a5[5][1] ;
 wire \CPU_Dmem_value_a5[5][20] ;
 wire \CPU_Dmem_value_a5[5][21] ;
 wire \CPU_Dmem_value_a5[5][22] ;
 wire \CPU_Dmem_value_a5[5][23] ;
 wire \CPU_Dmem_value_a5[5][24] ;
 wire \CPU_Dmem_value_a5[5][25] ;
 wire \CPU_Dmem_value_a5[5][26] ;
 wire \CPU_Dmem_value_a5[5][27] ;
 wire \CPU_Dmem_value_a5[5][28] ;
 wire \CPU_Dmem_value_a5[5][29] ;
 wire \CPU_Dmem_value_a5[5][2] ;
 wire \CPU_Dmem_value_a5[5][30] ;
 wire \CPU_Dmem_value_a5[5][31] ;
 wire \CPU_Dmem_value_a5[5][3] ;
 wire \CPU_Dmem_value_a5[5][4] ;
 wire \CPU_Dmem_value_a5[5][5] ;
 wire \CPU_Dmem_value_a5[5][6] ;
 wire \CPU_Dmem_value_a5[5][7] ;
 wire \CPU_Dmem_value_a5[5][8] ;
 wire \CPU_Dmem_value_a5[5][9] ;
 wire \CPU_Dmem_value_a5[6][0] ;
 wire \CPU_Dmem_value_a5[6][10] ;
 wire \CPU_Dmem_value_a5[6][11] ;
 wire \CPU_Dmem_value_a5[6][12] ;
 wire \CPU_Dmem_value_a5[6][13] ;
 wire \CPU_Dmem_value_a5[6][14] ;
 wire \CPU_Dmem_value_a5[6][15] ;
 wire \CPU_Dmem_value_a5[6][16] ;
 wire \CPU_Dmem_value_a5[6][17] ;
 wire \CPU_Dmem_value_a5[6][18] ;
 wire \CPU_Dmem_value_a5[6][19] ;
 wire \CPU_Dmem_value_a5[6][1] ;
 wire \CPU_Dmem_value_a5[6][20] ;
 wire \CPU_Dmem_value_a5[6][21] ;
 wire \CPU_Dmem_value_a5[6][22] ;
 wire \CPU_Dmem_value_a5[6][23] ;
 wire \CPU_Dmem_value_a5[6][24] ;
 wire \CPU_Dmem_value_a5[6][25] ;
 wire \CPU_Dmem_value_a5[6][26] ;
 wire \CPU_Dmem_value_a5[6][27] ;
 wire \CPU_Dmem_value_a5[6][28] ;
 wire \CPU_Dmem_value_a5[6][29] ;
 wire \CPU_Dmem_value_a5[6][2] ;
 wire \CPU_Dmem_value_a5[6][30] ;
 wire \CPU_Dmem_value_a5[6][31] ;
 wire \CPU_Dmem_value_a5[6][3] ;
 wire \CPU_Dmem_value_a5[6][4] ;
 wire \CPU_Dmem_value_a5[6][5] ;
 wire \CPU_Dmem_value_a5[6][6] ;
 wire \CPU_Dmem_value_a5[6][7] ;
 wire \CPU_Dmem_value_a5[6][8] ;
 wire \CPU_Dmem_value_a5[6][9] ;
 wire \CPU_Dmem_value_a5[7][0] ;
 wire \CPU_Dmem_value_a5[7][10] ;
 wire \CPU_Dmem_value_a5[7][11] ;
 wire \CPU_Dmem_value_a5[7][12] ;
 wire \CPU_Dmem_value_a5[7][13] ;
 wire \CPU_Dmem_value_a5[7][14] ;
 wire \CPU_Dmem_value_a5[7][15] ;
 wire \CPU_Dmem_value_a5[7][16] ;
 wire \CPU_Dmem_value_a5[7][17] ;
 wire \CPU_Dmem_value_a5[7][18] ;
 wire \CPU_Dmem_value_a5[7][19] ;
 wire \CPU_Dmem_value_a5[7][1] ;
 wire \CPU_Dmem_value_a5[7][20] ;
 wire \CPU_Dmem_value_a5[7][21] ;
 wire \CPU_Dmem_value_a5[7][22] ;
 wire \CPU_Dmem_value_a5[7][23] ;
 wire \CPU_Dmem_value_a5[7][24] ;
 wire \CPU_Dmem_value_a5[7][25] ;
 wire \CPU_Dmem_value_a5[7][26] ;
 wire \CPU_Dmem_value_a5[7][27] ;
 wire \CPU_Dmem_value_a5[7][28] ;
 wire \CPU_Dmem_value_a5[7][29] ;
 wire \CPU_Dmem_value_a5[7][2] ;
 wire \CPU_Dmem_value_a5[7][30] ;
 wire \CPU_Dmem_value_a5[7][31] ;
 wire \CPU_Dmem_value_a5[7][3] ;
 wire \CPU_Dmem_value_a5[7][4] ;
 wire \CPU_Dmem_value_a5[7][5] ;
 wire \CPU_Dmem_value_a5[7][6] ;
 wire \CPU_Dmem_value_a5[7][7] ;
 wire \CPU_Dmem_value_a5[7][8] ;
 wire \CPU_Dmem_value_a5[7][9] ;
 wire \CPU_Dmem_value_a5[8][0] ;
 wire \CPU_Dmem_value_a5[8][10] ;
 wire \CPU_Dmem_value_a5[8][11] ;
 wire \CPU_Dmem_value_a5[8][12] ;
 wire \CPU_Dmem_value_a5[8][13] ;
 wire \CPU_Dmem_value_a5[8][14] ;
 wire \CPU_Dmem_value_a5[8][15] ;
 wire \CPU_Dmem_value_a5[8][16] ;
 wire \CPU_Dmem_value_a5[8][17] ;
 wire \CPU_Dmem_value_a5[8][18] ;
 wire \CPU_Dmem_value_a5[8][19] ;
 wire \CPU_Dmem_value_a5[8][1] ;
 wire \CPU_Dmem_value_a5[8][20] ;
 wire \CPU_Dmem_value_a5[8][21] ;
 wire \CPU_Dmem_value_a5[8][22] ;
 wire \CPU_Dmem_value_a5[8][23] ;
 wire \CPU_Dmem_value_a5[8][24] ;
 wire \CPU_Dmem_value_a5[8][25] ;
 wire \CPU_Dmem_value_a5[8][26] ;
 wire \CPU_Dmem_value_a5[8][27] ;
 wire \CPU_Dmem_value_a5[8][28] ;
 wire \CPU_Dmem_value_a5[8][29] ;
 wire \CPU_Dmem_value_a5[8][2] ;
 wire \CPU_Dmem_value_a5[8][30] ;
 wire \CPU_Dmem_value_a5[8][31] ;
 wire \CPU_Dmem_value_a5[8][3] ;
 wire \CPU_Dmem_value_a5[8][4] ;
 wire \CPU_Dmem_value_a5[8][5] ;
 wire \CPU_Dmem_value_a5[8][6] ;
 wire \CPU_Dmem_value_a5[8][7] ;
 wire \CPU_Dmem_value_a5[8][8] ;
 wire \CPU_Dmem_value_a5[8][9] ;
 wire \CPU_Dmem_value_a5[9][0] ;
 wire \CPU_Dmem_value_a5[9][10] ;
 wire \CPU_Dmem_value_a5[9][11] ;
 wire \CPU_Dmem_value_a5[9][12] ;
 wire \CPU_Dmem_value_a5[9][13] ;
 wire \CPU_Dmem_value_a5[9][14] ;
 wire \CPU_Dmem_value_a5[9][15] ;
 wire \CPU_Dmem_value_a5[9][16] ;
 wire \CPU_Dmem_value_a5[9][17] ;
 wire \CPU_Dmem_value_a5[9][18] ;
 wire \CPU_Dmem_value_a5[9][19] ;
 wire \CPU_Dmem_value_a5[9][1] ;
 wire \CPU_Dmem_value_a5[9][20] ;
 wire \CPU_Dmem_value_a5[9][21] ;
 wire \CPU_Dmem_value_a5[9][22] ;
 wire \CPU_Dmem_value_a5[9][23] ;
 wire \CPU_Dmem_value_a5[9][24] ;
 wire \CPU_Dmem_value_a5[9][25] ;
 wire \CPU_Dmem_value_a5[9][26] ;
 wire \CPU_Dmem_value_a5[9][27] ;
 wire \CPU_Dmem_value_a5[9][28] ;
 wire \CPU_Dmem_value_a5[9][29] ;
 wire \CPU_Dmem_value_a5[9][2] ;
 wire \CPU_Dmem_value_a5[9][30] ;
 wire \CPU_Dmem_value_a5[9][31] ;
 wire \CPU_Dmem_value_a5[9][3] ;
 wire \CPU_Dmem_value_a5[9][4] ;
 wire \CPU_Dmem_value_a5[9][5] ;
 wire \CPU_Dmem_value_a5[9][6] ;
 wire \CPU_Dmem_value_a5[9][7] ;
 wire \CPU_Dmem_value_a5[9][8] ;
 wire \CPU_Dmem_value_a5[9][9] ;
 wire \CPU_Xreg_value_a4[0][0] ;
 wire \CPU_Xreg_value_a4[0][10] ;
 wire \CPU_Xreg_value_a4[0][11] ;
 wire \CPU_Xreg_value_a4[0][12] ;
 wire \CPU_Xreg_value_a4[0][13] ;
 wire \CPU_Xreg_value_a4[0][14] ;
 wire \CPU_Xreg_value_a4[0][15] ;
 wire \CPU_Xreg_value_a4[0][16] ;
 wire \CPU_Xreg_value_a4[0][17] ;
 wire \CPU_Xreg_value_a4[0][18] ;
 wire \CPU_Xreg_value_a4[0][19] ;
 wire \CPU_Xreg_value_a4[0][1] ;
 wire \CPU_Xreg_value_a4[0][20] ;
 wire \CPU_Xreg_value_a4[0][21] ;
 wire \CPU_Xreg_value_a4[0][22] ;
 wire \CPU_Xreg_value_a4[0][23] ;
 wire \CPU_Xreg_value_a4[0][24] ;
 wire \CPU_Xreg_value_a4[0][25] ;
 wire \CPU_Xreg_value_a4[0][26] ;
 wire \CPU_Xreg_value_a4[0][27] ;
 wire \CPU_Xreg_value_a4[0][28] ;
 wire \CPU_Xreg_value_a4[0][29] ;
 wire \CPU_Xreg_value_a4[0][2] ;
 wire \CPU_Xreg_value_a4[0][30] ;
 wire \CPU_Xreg_value_a4[0][31] ;
 wire \CPU_Xreg_value_a4[0][3] ;
 wire \CPU_Xreg_value_a4[0][4] ;
 wire \CPU_Xreg_value_a4[0][5] ;
 wire \CPU_Xreg_value_a4[0][6] ;
 wire \CPU_Xreg_value_a4[0][7] ;
 wire \CPU_Xreg_value_a4[0][8] ;
 wire \CPU_Xreg_value_a4[0][9] ;
 wire \CPU_Xreg_value_a4[10][0] ;
 wire \CPU_Xreg_value_a4[10][10] ;
 wire \CPU_Xreg_value_a4[10][11] ;
 wire \CPU_Xreg_value_a4[10][12] ;
 wire \CPU_Xreg_value_a4[10][13] ;
 wire \CPU_Xreg_value_a4[10][14] ;
 wire \CPU_Xreg_value_a4[10][15] ;
 wire \CPU_Xreg_value_a4[10][16] ;
 wire \CPU_Xreg_value_a4[10][17] ;
 wire \CPU_Xreg_value_a4[10][18] ;
 wire \CPU_Xreg_value_a4[10][19] ;
 wire \CPU_Xreg_value_a4[10][1] ;
 wire \CPU_Xreg_value_a4[10][20] ;
 wire \CPU_Xreg_value_a4[10][21] ;
 wire \CPU_Xreg_value_a4[10][22] ;
 wire \CPU_Xreg_value_a4[10][23] ;
 wire \CPU_Xreg_value_a4[10][24] ;
 wire \CPU_Xreg_value_a4[10][25] ;
 wire \CPU_Xreg_value_a4[10][26] ;
 wire \CPU_Xreg_value_a4[10][27] ;
 wire \CPU_Xreg_value_a4[10][28] ;
 wire \CPU_Xreg_value_a4[10][29] ;
 wire \CPU_Xreg_value_a4[10][2] ;
 wire \CPU_Xreg_value_a4[10][30] ;
 wire \CPU_Xreg_value_a4[10][31] ;
 wire \CPU_Xreg_value_a4[10][3] ;
 wire \CPU_Xreg_value_a4[10][4] ;
 wire \CPU_Xreg_value_a4[10][5] ;
 wire \CPU_Xreg_value_a4[10][6] ;
 wire \CPU_Xreg_value_a4[10][7] ;
 wire \CPU_Xreg_value_a4[10][8] ;
 wire \CPU_Xreg_value_a4[10][9] ;
 wire \CPU_Xreg_value_a4[11][0] ;
 wire \CPU_Xreg_value_a4[11][10] ;
 wire \CPU_Xreg_value_a4[11][11] ;
 wire \CPU_Xreg_value_a4[11][12] ;
 wire \CPU_Xreg_value_a4[11][13] ;
 wire \CPU_Xreg_value_a4[11][14] ;
 wire \CPU_Xreg_value_a4[11][15] ;
 wire \CPU_Xreg_value_a4[11][16] ;
 wire \CPU_Xreg_value_a4[11][17] ;
 wire \CPU_Xreg_value_a4[11][18] ;
 wire \CPU_Xreg_value_a4[11][19] ;
 wire \CPU_Xreg_value_a4[11][1] ;
 wire \CPU_Xreg_value_a4[11][20] ;
 wire \CPU_Xreg_value_a4[11][21] ;
 wire \CPU_Xreg_value_a4[11][22] ;
 wire \CPU_Xreg_value_a4[11][23] ;
 wire \CPU_Xreg_value_a4[11][24] ;
 wire \CPU_Xreg_value_a4[11][25] ;
 wire \CPU_Xreg_value_a4[11][26] ;
 wire \CPU_Xreg_value_a4[11][27] ;
 wire \CPU_Xreg_value_a4[11][28] ;
 wire \CPU_Xreg_value_a4[11][29] ;
 wire \CPU_Xreg_value_a4[11][2] ;
 wire \CPU_Xreg_value_a4[11][30] ;
 wire \CPU_Xreg_value_a4[11][31] ;
 wire \CPU_Xreg_value_a4[11][3] ;
 wire \CPU_Xreg_value_a4[11][4] ;
 wire \CPU_Xreg_value_a4[11][5] ;
 wire \CPU_Xreg_value_a4[11][6] ;
 wire \CPU_Xreg_value_a4[11][7] ;
 wire \CPU_Xreg_value_a4[11][8] ;
 wire \CPU_Xreg_value_a4[11][9] ;
 wire \CPU_Xreg_value_a4[12][0] ;
 wire \CPU_Xreg_value_a4[12][10] ;
 wire \CPU_Xreg_value_a4[12][11] ;
 wire \CPU_Xreg_value_a4[12][12] ;
 wire \CPU_Xreg_value_a4[12][13] ;
 wire \CPU_Xreg_value_a4[12][14] ;
 wire \CPU_Xreg_value_a4[12][15] ;
 wire \CPU_Xreg_value_a4[12][16] ;
 wire \CPU_Xreg_value_a4[12][17] ;
 wire \CPU_Xreg_value_a4[12][18] ;
 wire \CPU_Xreg_value_a4[12][19] ;
 wire \CPU_Xreg_value_a4[12][1] ;
 wire \CPU_Xreg_value_a4[12][20] ;
 wire \CPU_Xreg_value_a4[12][21] ;
 wire \CPU_Xreg_value_a4[12][22] ;
 wire \CPU_Xreg_value_a4[12][23] ;
 wire \CPU_Xreg_value_a4[12][24] ;
 wire \CPU_Xreg_value_a4[12][25] ;
 wire \CPU_Xreg_value_a4[12][26] ;
 wire \CPU_Xreg_value_a4[12][27] ;
 wire \CPU_Xreg_value_a4[12][28] ;
 wire \CPU_Xreg_value_a4[12][29] ;
 wire \CPU_Xreg_value_a4[12][2] ;
 wire \CPU_Xreg_value_a4[12][30] ;
 wire \CPU_Xreg_value_a4[12][31] ;
 wire \CPU_Xreg_value_a4[12][3] ;
 wire \CPU_Xreg_value_a4[12][4] ;
 wire \CPU_Xreg_value_a4[12][5] ;
 wire \CPU_Xreg_value_a4[12][6] ;
 wire \CPU_Xreg_value_a4[12][7] ;
 wire \CPU_Xreg_value_a4[12][8] ;
 wire \CPU_Xreg_value_a4[12][9] ;
 wire \CPU_Xreg_value_a4[13][0] ;
 wire \CPU_Xreg_value_a4[13][10] ;
 wire \CPU_Xreg_value_a4[13][11] ;
 wire \CPU_Xreg_value_a4[13][12] ;
 wire \CPU_Xreg_value_a4[13][13] ;
 wire \CPU_Xreg_value_a4[13][14] ;
 wire \CPU_Xreg_value_a4[13][15] ;
 wire \CPU_Xreg_value_a4[13][16] ;
 wire \CPU_Xreg_value_a4[13][17] ;
 wire \CPU_Xreg_value_a4[13][18] ;
 wire \CPU_Xreg_value_a4[13][19] ;
 wire \CPU_Xreg_value_a4[13][1] ;
 wire \CPU_Xreg_value_a4[13][20] ;
 wire \CPU_Xreg_value_a4[13][21] ;
 wire \CPU_Xreg_value_a4[13][22] ;
 wire \CPU_Xreg_value_a4[13][23] ;
 wire \CPU_Xreg_value_a4[13][24] ;
 wire \CPU_Xreg_value_a4[13][25] ;
 wire \CPU_Xreg_value_a4[13][26] ;
 wire \CPU_Xreg_value_a4[13][27] ;
 wire \CPU_Xreg_value_a4[13][28] ;
 wire \CPU_Xreg_value_a4[13][29] ;
 wire \CPU_Xreg_value_a4[13][2] ;
 wire \CPU_Xreg_value_a4[13][30] ;
 wire \CPU_Xreg_value_a4[13][31] ;
 wire \CPU_Xreg_value_a4[13][3] ;
 wire \CPU_Xreg_value_a4[13][4] ;
 wire \CPU_Xreg_value_a4[13][5] ;
 wire \CPU_Xreg_value_a4[13][6] ;
 wire \CPU_Xreg_value_a4[13][7] ;
 wire \CPU_Xreg_value_a4[13][8] ;
 wire \CPU_Xreg_value_a4[13][9] ;
 wire \CPU_Xreg_value_a4[14][0] ;
 wire \CPU_Xreg_value_a4[14][10] ;
 wire \CPU_Xreg_value_a4[14][11] ;
 wire \CPU_Xreg_value_a4[14][12] ;
 wire \CPU_Xreg_value_a4[14][13] ;
 wire \CPU_Xreg_value_a4[14][14] ;
 wire \CPU_Xreg_value_a4[14][15] ;
 wire \CPU_Xreg_value_a4[14][16] ;
 wire \CPU_Xreg_value_a4[14][17] ;
 wire \CPU_Xreg_value_a4[14][18] ;
 wire \CPU_Xreg_value_a4[14][19] ;
 wire \CPU_Xreg_value_a4[14][1] ;
 wire \CPU_Xreg_value_a4[14][20] ;
 wire \CPU_Xreg_value_a4[14][21] ;
 wire \CPU_Xreg_value_a4[14][22] ;
 wire \CPU_Xreg_value_a4[14][23] ;
 wire \CPU_Xreg_value_a4[14][24] ;
 wire \CPU_Xreg_value_a4[14][25] ;
 wire \CPU_Xreg_value_a4[14][26] ;
 wire \CPU_Xreg_value_a4[14][27] ;
 wire \CPU_Xreg_value_a4[14][28] ;
 wire \CPU_Xreg_value_a4[14][29] ;
 wire \CPU_Xreg_value_a4[14][2] ;
 wire \CPU_Xreg_value_a4[14][30] ;
 wire \CPU_Xreg_value_a4[14][31] ;
 wire \CPU_Xreg_value_a4[14][3] ;
 wire \CPU_Xreg_value_a4[14][4] ;
 wire \CPU_Xreg_value_a4[14][5] ;
 wire \CPU_Xreg_value_a4[14][6] ;
 wire \CPU_Xreg_value_a4[14][7] ;
 wire \CPU_Xreg_value_a4[14][8] ;
 wire \CPU_Xreg_value_a4[14][9] ;
 wire \CPU_Xreg_value_a4[15][0] ;
 wire \CPU_Xreg_value_a4[15][10] ;
 wire \CPU_Xreg_value_a4[15][11] ;
 wire \CPU_Xreg_value_a4[15][12] ;
 wire \CPU_Xreg_value_a4[15][13] ;
 wire \CPU_Xreg_value_a4[15][14] ;
 wire \CPU_Xreg_value_a4[15][15] ;
 wire \CPU_Xreg_value_a4[15][16] ;
 wire \CPU_Xreg_value_a4[15][17] ;
 wire \CPU_Xreg_value_a4[15][18] ;
 wire \CPU_Xreg_value_a4[15][19] ;
 wire \CPU_Xreg_value_a4[15][1] ;
 wire \CPU_Xreg_value_a4[15][20] ;
 wire \CPU_Xreg_value_a4[15][21] ;
 wire \CPU_Xreg_value_a4[15][22] ;
 wire \CPU_Xreg_value_a4[15][23] ;
 wire \CPU_Xreg_value_a4[15][24] ;
 wire \CPU_Xreg_value_a4[15][25] ;
 wire \CPU_Xreg_value_a4[15][26] ;
 wire \CPU_Xreg_value_a4[15][27] ;
 wire \CPU_Xreg_value_a4[15][28] ;
 wire \CPU_Xreg_value_a4[15][29] ;
 wire \CPU_Xreg_value_a4[15][2] ;
 wire \CPU_Xreg_value_a4[15][30] ;
 wire \CPU_Xreg_value_a4[15][31] ;
 wire \CPU_Xreg_value_a4[15][3] ;
 wire \CPU_Xreg_value_a4[15][4] ;
 wire \CPU_Xreg_value_a4[15][5] ;
 wire \CPU_Xreg_value_a4[15][6] ;
 wire \CPU_Xreg_value_a4[15][7] ;
 wire \CPU_Xreg_value_a4[15][8] ;
 wire \CPU_Xreg_value_a4[15][9] ;
 wire \CPU_Xreg_value_a4[1][0] ;
 wire \CPU_Xreg_value_a4[1][10] ;
 wire \CPU_Xreg_value_a4[1][11] ;
 wire \CPU_Xreg_value_a4[1][12] ;
 wire \CPU_Xreg_value_a4[1][13] ;
 wire \CPU_Xreg_value_a4[1][14] ;
 wire \CPU_Xreg_value_a4[1][15] ;
 wire \CPU_Xreg_value_a4[1][16] ;
 wire \CPU_Xreg_value_a4[1][17] ;
 wire \CPU_Xreg_value_a4[1][18] ;
 wire \CPU_Xreg_value_a4[1][19] ;
 wire \CPU_Xreg_value_a4[1][1] ;
 wire \CPU_Xreg_value_a4[1][20] ;
 wire \CPU_Xreg_value_a4[1][21] ;
 wire \CPU_Xreg_value_a4[1][22] ;
 wire \CPU_Xreg_value_a4[1][23] ;
 wire \CPU_Xreg_value_a4[1][24] ;
 wire \CPU_Xreg_value_a4[1][25] ;
 wire \CPU_Xreg_value_a4[1][26] ;
 wire \CPU_Xreg_value_a4[1][27] ;
 wire \CPU_Xreg_value_a4[1][28] ;
 wire \CPU_Xreg_value_a4[1][29] ;
 wire \CPU_Xreg_value_a4[1][2] ;
 wire \CPU_Xreg_value_a4[1][30] ;
 wire \CPU_Xreg_value_a4[1][31] ;
 wire \CPU_Xreg_value_a4[1][3] ;
 wire \CPU_Xreg_value_a4[1][4] ;
 wire \CPU_Xreg_value_a4[1][5] ;
 wire \CPU_Xreg_value_a4[1][6] ;
 wire \CPU_Xreg_value_a4[1][7] ;
 wire \CPU_Xreg_value_a4[1][8] ;
 wire \CPU_Xreg_value_a4[1][9] ;
 wire \CPU_Xreg_value_a4[2][0] ;
 wire \CPU_Xreg_value_a4[2][10] ;
 wire \CPU_Xreg_value_a4[2][11] ;
 wire \CPU_Xreg_value_a4[2][12] ;
 wire \CPU_Xreg_value_a4[2][13] ;
 wire \CPU_Xreg_value_a4[2][14] ;
 wire \CPU_Xreg_value_a4[2][15] ;
 wire \CPU_Xreg_value_a4[2][16] ;
 wire \CPU_Xreg_value_a4[2][17] ;
 wire \CPU_Xreg_value_a4[2][18] ;
 wire \CPU_Xreg_value_a4[2][19] ;
 wire \CPU_Xreg_value_a4[2][1] ;
 wire \CPU_Xreg_value_a4[2][20] ;
 wire \CPU_Xreg_value_a4[2][21] ;
 wire \CPU_Xreg_value_a4[2][22] ;
 wire \CPU_Xreg_value_a4[2][23] ;
 wire \CPU_Xreg_value_a4[2][24] ;
 wire \CPU_Xreg_value_a4[2][25] ;
 wire \CPU_Xreg_value_a4[2][26] ;
 wire \CPU_Xreg_value_a4[2][27] ;
 wire \CPU_Xreg_value_a4[2][28] ;
 wire \CPU_Xreg_value_a4[2][29] ;
 wire \CPU_Xreg_value_a4[2][2] ;
 wire \CPU_Xreg_value_a4[2][30] ;
 wire \CPU_Xreg_value_a4[2][31] ;
 wire \CPU_Xreg_value_a4[2][3] ;
 wire \CPU_Xreg_value_a4[2][4] ;
 wire \CPU_Xreg_value_a4[2][5] ;
 wire \CPU_Xreg_value_a4[2][6] ;
 wire \CPU_Xreg_value_a4[2][7] ;
 wire \CPU_Xreg_value_a4[2][8] ;
 wire \CPU_Xreg_value_a4[2][9] ;
 wire \CPU_Xreg_value_a4[3][0] ;
 wire \CPU_Xreg_value_a4[3][10] ;
 wire \CPU_Xreg_value_a4[3][11] ;
 wire \CPU_Xreg_value_a4[3][12] ;
 wire \CPU_Xreg_value_a4[3][13] ;
 wire \CPU_Xreg_value_a4[3][14] ;
 wire \CPU_Xreg_value_a4[3][15] ;
 wire \CPU_Xreg_value_a4[3][16] ;
 wire \CPU_Xreg_value_a4[3][17] ;
 wire \CPU_Xreg_value_a4[3][18] ;
 wire \CPU_Xreg_value_a4[3][19] ;
 wire \CPU_Xreg_value_a4[3][1] ;
 wire \CPU_Xreg_value_a4[3][20] ;
 wire \CPU_Xreg_value_a4[3][21] ;
 wire \CPU_Xreg_value_a4[3][22] ;
 wire \CPU_Xreg_value_a4[3][23] ;
 wire \CPU_Xreg_value_a4[3][24] ;
 wire \CPU_Xreg_value_a4[3][25] ;
 wire \CPU_Xreg_value_a4[3][26] ;
 wire \CPU_Xreg_value_a4[3][27] ;
 wire \CPU_Xreg_value_a4[3][28] ;
 wire \CPU_Xreg_value_a4[3][29] ;
 wire \CPU_Xreg_value_a4[3][2] ;
 wire \CPU_Xreg_value_a4[3][30] ;
 wire \CPU_Xreg_value_a4[3][31] ;
 wire \CPU_Xreg_value_a4[3][3] ;
 wire \CPU_Xreg_value_a4[3][4] ;
 wire \CPU_Xreg_value_a4[3][5] ;
 wire \CPU_Xreg_value_a4[3][6] ;
 wire \CPU_Xreg_value_a4[3][7] ;
 wire \CPU_Xreg_value_a4[3][8] ;
 wire \CPU_Xreg_value_a4[3][9] ;
 wire \CPU_Xreg_value_a4[4][0] ;
 wire \CPU_Xreg_value_a4[4][10] ;
 wire \CPU_Xreg_value_a4[4][11] ;
 wire \CPU_Xreg_value_a4[4][12] ;
 wire \CPU_Xreg_value_a4[4][13] ;
 wire \CPU_Xreg_value_a4[4][14] ;
 wire \CPU_Xreg_value_a4[4][15] ;
 wire \CPU_Xreg_value_a4[4][16] ;
 wire \CPU_Xreg_value_a4[4][17] ;
 wire \CPU_Xreg_value_a4[4][18] ;
 wire \CPU_Xreg_value_a4[4][19] ;
 wire \CPU_Xreg_value_a4[4][1] ;
 wire \CPU_Xreg_value_a4[4][20] ;
 wire \CPU_Xreg_value_a4[4][21] ;
 wire \CPU_Xreg_value_a4[4][22] ;
 wire \CPU_Xreg_value_a4[4][23] ;
 wire \CPU_Xreg_value_a4[4][24] ;
 wire \CPU_Xreg_value_a4[4][25] ;
 wire \CPU_Xreg_value_a4[4][26] ;
 wire \CPU_Xreg_value_a4[4][27] ;
 wire \CPU_Xreg_value_a4[4][28] ;
 wire \CPU_Xreg_value_a4[4][29] ;
 wire \CPU_Xreg_value_a4[4][2] ;
 wire \CPU_Xreg_value_a4[4][30] ;
 wire \CPU_Xreg_value_a4[4][31] ;
 wire \CPU_Xreg_value_a4[4][3] ;
 wire \CPU_Xreg_value_a4[4][4] ;
 wire \CPU_Xreg_value_a4[4][5] ;
 wire \CPU_Xreg_value_a4[4][6] ;
 wire \CPU_Xreg_value_a4[4][7] ;
 wire \CPU_Xreg_value_a4[4][8] ;
 wire \CPU_Xreg_value_a4[4][9] ;
 wire \CPU_Xreg_value_a4[5][0] ;
 wire \CPU_Xreg_value_a4[5][10] ;
 wire \CPU_Xreg_value_a4[5][11] ;
 wire \CPU_Xreg_value_a4[5][12] ;
 wire \CPU_Xreg_value_a4[5][13] ;
 wire \CPU_Xreg_value_a4[5][14] ;
 wire \CPU_Xreg_value_a4[5][15] ;
 wire \CPU_Xreg_value_a4[5][16] ;
 wire \CPU_Xreg_value_a4[5][17] ;
 wire \CPU_Xreg_value_a4[5][18] ;
 wire \CPU_Xreg_value_a4[5][19] ;
 wire \CPU_Xreg_value_a4[5][1] ;
 wire \CPU_Xreg_value_a4[5][20] ;
 wire \CPU_Xreg_value_a4[5][21] ;
 wire \CPU_Xreg_value_a4[5][22] ;
 wire \CPU_Xreg_value_a4[5][23] ;
 wire \CPU_Xreg_value_a4[5][24] ;
 wire \CPU_Xreg_value_a4[5][25] ;
 wire \CPU_Xreg_value_a4[5][26] ;
 wire \CPU_Xreg_value_a4[5][27] ;
 wire \CPU_Xreg_value_a4[5][28] ;
 wire \CPU_Xreg_value_a4[5][29] ;
 wire \CPU_Xreg_value_a4[5][2] ;
 wire \CPU_Xreg_value_a4[5][30] ;
 wire \CPU_Xreg_value_a4[5][31] ;
 wire \CPU_Xreg_value_a4[5][3] ;
 wire \CPU_Xreg_value_a4[5][4] ;
 wire \CPU_Xreg_value_a4[5][5] ;
 wire \CPU_Xreg_value_a4[5][6] ;
 wire \CPU_Xreg_value_a4[5][7] ;
 wire \CPU_Xreg_value_a4[5][8] ;
 wire \CPU_Xreg_value_a4[5][9] ;
 wire \CPU_Xreg_value_a4[6][0] ;
 wire \CPU_Xreg_value_a4[6][10] ;
 wire \CPU_Xreg_value_a4[6][11] ;
 wire \CPU_Xreg_value_a4[6][12] ;
 wire \CPU_Xreg_value_a4[6][13] ;
 wire \CPU_Xreg_value_a4[6][14] ;
 wire \CPU_Xreg_value_a4[6][15] ;
 wire \CPU_Xreg_value_a4[6][16] ;
 wire \CPU_Xreg_value_a4[6][17] ;
 wire \CPU_Xreg_value_a4[6][18] ;
 wire \CPU_Xreg_value_a4[6][19] ;
 wire \CPU_Xreg_value_a4[6][1] ;
 wire \CPU_Xreg_value_a4[6][20] ;
 wire \CPU_Xreg_value_a4[6][21] ;
 wire \CPU_Xreg_value_a4[6][22] ;
 wire \CPU_Xreg_value_a4[6][23] ;
 wire \CPU_Xreg_value_a4[6][24] ;
 wire \CPU_Xreg_value_a4[6][25] ;
 wire \CPU_Xreg_value_a4[6][26] ;
 wire \CPU_Xreg_value_a4[6][27] ;
 wire \CPU_Xreg_value_a4[6][28] ;
 wire \CPU_Xreg_value_a4[6][29] ;
 wire \CPU_Xreg_value_a4[6][2] ;
 wire \CPU_Xreg_value_a4[6][30] ;
 wire \CPU_Xreg_value_a4[6][31] ;
 wire \CPU_Xreg_value_a4[6][3] ;
 wire \CPU_Xreg_value_a4[6][4] ;
 wire \CPU_Xreg_value_a4[6][5] ;
 wire \CPU_Xreg_value_a4[6][6] ;
 wire \CPU_Xreg_value_a4[6][7] ;
 wire \CPU_Xreg_value_a4[6][8] ;
 wire \CPU_Xreg_value_a4[6][9] ;
 wire \CPU_Xreg_value_a4[7][0] ;
 wire \CPU_Xreg_value_a4[7][10] ;
 wire \CPU_Xreg_value_a4[7][11] ;
 wire \CPU_Xreg_value_a4[7][12] ;
 wire \CPU_Xreg_value_a4[7][13] ;
 wire \CPU_Xreg_value_a4[7][14] ;
 wire \CPU_Xreg_value_a4[7][15] ;
 wire \CPU_Xreg_value_a4[7][16] ;
 wire \CPU_Xreg_value_a4[7][17] ;
 wire \CPU_Xreg_value_a4[7][18] ;
 wire \CPU_Xreg_value_a4[7][19] ;
 wire \CPU_Xreg_value_a4[7][1] ;
 wire \CPU_Xreg_value_a4[7][20] ;
 wire \CPU_Xreg_value_a4[7][21] ;
 wire \CPU_Xreg_value_a4[7][22] ;
 wire \CPU_Xreg_value_a4[7][23] ;
 wire \CPU_Xreg_value_a4[7][24] ;
 wire \CPU_Xreg_value_a4[7][25] ;
 wire \CPU_Xreg_value_a4[7][26] ;
 wire \CPU_Xreg_value_a4[7][27] ;
 wire \CPU_Xreg_value_a4[7][28] ;
 wire \CPU_Xreg_value_a4[7][29] ;
 wire \CPU_Xreg_value_a4[7][2] ;
 wire \CPU_Xreg_value_a4[7][30] ;
 wire \CPU_Xreg_value_a4[7][31] ;
 wire \CPU_Xreg_value_a4[7][3] ;
 wire \CPU_Xreg_value_a4[7][4] ;
 wire \CPU_Xreg_value_a4[7][5] ;
 wire \CPU_Xreg_value_a4[7][6] ;
 wire \CPU_Xreg_value_a4[7][7] ;
 wire \CPU_Xreg_value_a4[7][8] ;
 wire \CPU_Xreg_value_a4[7][9] ;
 wire \CPU_Xreg_value_a4[8][0] ;
 wire \CPU_Xreg_value_a4[8][10] ;
 wire \CPU_Xreg_value_a4[8][11] ;
 wire \CPU_Xreg_value_a4[8][12] ;
 wire \CPU_Xreg_value_a4[8][13] ;
 wire \CPU_Xreg_value_a4[8][14] ;
 wire \CPU_Xreg_value_a4[8][15] ;
 wire \CPU_Xreg_value_a4[8][16] ;
 wire \CPU_Xreg_value_a4[8][17] ;
 wire \CPU_Xreg_value_a4[8][18] ;
 wire \CPU_Xreg_value_a4[8][19] ;
 wire \CPU_Xreg_value_a4[8][1] ;
 wire \CPU_Xreg_value_a4[8][20] ;
 wire \CPU_Xreg_value_a4[8][21] ;
 wire \CPU_Xreg_value_a4[8][22] ;
 wire \CPU_Xreg_value_a4[8][23] ;
 wire \CPU_Xreg_value_a4[8][24] ;
 wire \CPU_Xreg_value_a4[8][25] ;
 wire \CPU_Xreg_value_a4[8][26] ;
 wire \CPU_Xreg_value_a4[8][27] ;
 wire \CPU_Xreg_value_a4[8][28] ;
 wire \CPU_Xreg_value_a4[8][29] ;
 wire \CPU_Xreg_value_a4[8][2] ;
 wire \CPU_Xreg_value_a4[8][30] ;
 wire \CPU_Xreg_value_a4[8][31] ;
 wire \CPU_Xreg_value_a4[8][3] ;
 wire \CPU_Xreg_value_a4[8][4] ;
 wire \CPU_Xreg_value_a4[8][5] ;
 wire \CPU_Xreg_value_a4[8][6] ;
 wire \CPU_Xreg_value_a4[8][7] ;
 wire \CPU_Xreg_value_a4[8][8] ;
 wire \CPU_Xreg_value_a4[8][9] ;
 wire \CPU_Xreg_value_a4[9][0] ;
 wire \CPU_Xreg_value_a4[9][10] ;
 wire \CPU_Xreg_value_a4[9][11] ;
 wire \CPU_Xreg_value_a4[9][12] ;
 wire \CPU_Xreg_value_a4[9][13] ;
 wire \CPU_Xreg_value_a4[9][14] ;
 wire \CPU_Xreg_value_a4[9][15] ;
 wire \CPU_Xreg_value_a4[9][16] ;
 wire \CPU_Xreg_value_a4[9][17] ;
 wire \CPU_Xreg_value_a4[9][18] ;
 wire \CPU_Xreg_value_a4[9][19] ;
 wire \CPU_Xreg_value_a4[9][1] ;
 wire \CPU_Xreg_value_a4[9][20] ;
 wire \CPU_Xreg_value_a4[9][21] ;
 wire \CPU_Xreg_value_a4[9][22] ;
 wire \CPU_Xreg_value_a4[9][23] ;
 wire \CPU_Xreg_value_a4[9][24] ;
 wire \CPU_Xreg_value_a4[9][25] ;
 wire \CPU_Xreg_value_a4[9][26] ;
 wire \CPU_Xreg_value_a4[9][27] ;
 wire \CPU_Xreg_value_a4[9][28] ;
 wire \CPU_Xreg_value_a4[9][29] ;
 wire \CPU_Xreg_value_a4[9][2] ;
 wire \CPU_Xreg_value_a4[9][30] ;
 wire \CPU_Xreg_value_a4[9][31] ;
 wire \CPU_Xreg_value_a4[9][3] ;
 wire \CPU_Xreg_value_a4[9][4] ;
 wire \CPU_Xreg_value_a4[9][5] ;
 wire \CPU_Xreg_value_a4[9][6] ;
 wire \CPU_Xreg_value_a4[9][7] ;
 wire \CPU_Xreg_value_a4[9][8] ;
 wire \CPU_Xreg_value_a4[9][9] ;
 wire \CPU_Xreg_value_a5[14][0] ;
 wire \CPU_Xreg_value_a5[14][1] ;
 wire \CPU_Xreg_value_a5[14][2] ;
 wire \CPU_Xreg_value_a5[14][3] ;
 wire \CPU_Xreg_value_a5[14][4] ;
 wire \CPU_Xreg_value_a5[14][5] ;
 wire \CPU_Xreg_value_a5[14][6] ;
 wire \CPU_Xreg_value_a5[14][7] ;
 wire \CPU_Xreg_value_a5[14][8] ;
 wire \CPU_Xreg_value_a5[14][9] ;
 wire \CPU_br_tgt_pc_a2[0] ;
 wire \CPU_br_tgt_pc_a2[1] ;
 wire \CPU_br_tgt_pc_a2[2] ;
 wire \CPU_br_tgt_pc_a2[3] ;
 wire \CPU_br_tgt_pc_a2[4] ;
 wire \CPU_br_tgt_pc_a2[5] ;
 wire \CPU_br_tgt_pc_a3[0] ;
 wire \CPU_br_tgt_pc_a3[1] ;
 wire \CPU_br_tgt_pc_a3[2] ;
 wire \CPU_br_tgt_pc_a3[3] ;
 wire \CPU_br_tgt_pc_a3[4] ;
 wire \CPU_br_tgt_pc_a3[5] ;
 wire \CPU_dec_bits_a1[10] ;
 wire \CPU_dmem_addr_a4[0] ;
 wire \CPU_dmem_addr_a4[1] ;
 wire \CPU_dmem_addr_a4[2] ;
 wire \CPU_dmem_addr_a4[3] ;
 wire \CPU_dmem_rd_data_a5[0] ;
 wire \CPU_dmem_rd_data_a5[10] ;
 wire \CPU_dmem_rd_data_a5[11] ;
 wire \CPU_dmem_rd_data_a5[12] ;
 wire \CPU_dmem_rd_data_a5[13] ;
 wire \CPU_dmem_rd_data_a5[14] ;
 wire \CPU_dmem_rd_data_a5[15] ;
 wire \CPU_dmem_rd_data_a5[16] ;
 wire \CPU_dmem_rd_data_a5[17] ;
 wire \CPU_dmem_rd_data_a5[18] ;
 wire \CPU_dmem_rd_data_a5[19] ;
 wire \CPU_dmem_rd_data_a5[1] ;
 wire \CPU_dmem_rd_data_a5[20] ;
 wire \CPU_dmem_rd_data_a5[21] ;
 wire \CPU_dmem_rd_data_a5[22] ;
 wire \CPU_dmem_rd_data_a5[23] ;
 wire \CPU_dmem_rd_data_a5[24] ;
 wire \CPU_dmem_rd_data_a5[25] ;
 wire \CPU_dmem_rd_data_a5[26] ;
 wire \CPU_dmem_rd_data_a5[27] ;
 wire \CPU_dmem_rd_data_a5[28] ;
 wire \CPU_dmem_rd_data_a5[29] ;
 wire \CPU_dmem_rd_data_a5[2] ;
 wire \CPU_dmem_rd_data_a5[30] ;
 wire \CPU_dmem_rd_data_a5[31] ;
 wire \CPU_dmem_rd_data_a5[3] ;
 wire \CPU_dmem_rd_data_a5[4] ;
 wire \CPU_dmem_rd_data_a5[5] ;
 wire \CPU_dmem_rd_data_a5[6] ;
 wire \CPU_dmem_rd_data_a5[7] ;
 wire \CPU_dmem_rd_data_a5[8] ;
 wire \CPU_dmem_rd_data_a5[9] ;
 wire CPU_dmem_rd_en_a4;
 wire \CPU_dmem_wr_data_a4[0] ;
 wire \CPU_dmem_wr_data_a4[10] ;
 wire \CPU_dmem_wr_data_a4[11] ;
 wire \CPU_dmem_wr_data_a4[12] ;
 wire \CPU_dmem_wr_data_a4[13] ;
 wire \CPU_dmem_wr_data_a4[14] ;
 wire \CPU_dmem_wr_data_a4[15] ;
 wire \CPU_dmem_wr_data_a4[16] ;
 wire \CPU_dmem_wr_data_a4[17] ;
 wire \CPU_dmem_wr_data_a4[18] ;
 wire \CPU_dmem_wr_data_a4[19] ;
 wire \CPU_dmem_wr_data_a4[1] ;
 wire \CPU_dmem_wr_data_a4[20] ;
 wire \CPU_dmem_wr_data_a4[21] ;
 wire \CPU_dmem_wr_data_a4[22] ;
 wire \CPU_dmem_wr_data_a4[23] ;
 wire \CPU_dmem_wr_data_a4[24] ;
 wire \CPU_dmem_wr_data_a4[25] ;
 wire \CPU_dmem_wr_data_a4[26] ;
 wire \CPU_dmem_wr_data_a4[27] ;
 wire \CPU_dmem_wr_data_a4[28] ;
 wire \CPU_dmem_wr_data_a4[29] ;
 wire \CPU_dmem_wr_data_a4[2] ;
 wire \CPU_dmem_wr_data_a4[30] ;
 wire \CPU_dmem_wr_data_a4[31] ;
 wire \CPU_dmem_wr_data_a4[3] ;
 wire \CPU_dmem_wr_data_a4[4] ;
 wire \CPU_dmem_wr_data_a4[5] ;
 wire \CPU_dmem_wr_data_a4[6] ;
 wire \CPU_dmem_wr_data_a4[7] ;
 wire \CPU_dmem_wr_data_a4[8] ;
 wire \CPU_dmem_wr_data_a4[9] ;
 wire \CPU_imem_rd_addr_a1[0] ;
 wire \CPU_imem_rd_addr_a1[1] ;
 wire \CPU_imem_rd_addr_a1[2] ;
 wire \CPU_imem_rd_addr_a1[3] ;
 wire \CPU_imem_rd_data_a1[10] ;
 wire \CPU_imem_rd_data_a1[20] ;
 wire \CPU_imem_rd_data_a1[21] ;
 wire \CPU_imem_rd_data_a1[22] ;
 wire \CPU_imem_rd_data_a1[23] ;
 wire \CPU_imem_rd_data_a1[7] ;
 wire \CPU_imem_rd_data_a1[8] ;
 wire \CPU_imem_rd_data_a1[9] ;
 wire \CPU_imm_a1[0] ;
 wire \CPU_imm_a1[10] ;
 wire \CPU_imm_a1[11] ;
 wire \CPU_imm_a1[1] ;
 wire \CPU_imm_a1[2] ;
 wire \CPU_imm_a1[3] ;
 wire \CPU_imm_a2[0] ;
 wire \CPU_imm_a2[10] ;
 wire \CPU_imm_a2[11] ;
 wire \CPU_imm_a2[1] ;
 wire \CPU_imm_a2[2] ;
 wire \CPU_imm_a2[3] ;
 wire \CPU_imm_a2[4] ;
 wire \CPU_imm_a3[0] ;
 wire \CPU_imm_a3[10] ;
 wire \CPU_imm_a3[11] ;
 wire \CPU_imm_a3[1] ;
 wire \CPU_imm_a3[2] ;
 wire \CPU_imm_a3[3] ;
 wire \CPU_imm_a3[4] ;
 wire \CPU_inc_pc_a1[0] ;
 wire \CPU_inc_pc_a1[1] ;
 wire \CPU_inc_pc_a1[2] ;
 wire \CPU_inc_pc_a1[3] ;
 wire \CPU_inc_pc_a1[4] ;
 wire \CPU_inc_pc_a1[5] ;
 wire \CPU_inc_pc_a2[0] ;
 wire \CPU_inc_pc_a2[1] ;
 wire \CPU_inc_pc_a2[2] ;
 wire \CPU_inc_pc_a2[3] ;
 wire \CPU_inc_pc_a2[4] ;
 wire \CPU_inc_pc_a2[5] ;
 wire \CPU_inc_pc_a3[0] ;
 wire \CPU_inc_pc_a3[1] ;
 wire \CPU_inc_pc_a3[2] ;
 wire \CPU_inc_pc_a3[3] ;
 wire \CPU_inc_pc_a3[4] ;
 wire \CPU_inc_pc_a3[5] ;
 wire CPU_is_add_a1;
 wire CPU_is_add_a2;
 wire CPU_is_add_a3;
 wire CPU_is_addi_a1;
 wire CPU_is_addi_a2;
 wire CPU_is_addi_a3;
 wire CPU_is_blt_a1;
 wire CPU_is_blt_a2;
 wire CPU_is_blt_a3;
 wire CPU_is_bltu_a2;
 wire CPU_is_bltu_a3;
 wire CPU_is_load_a1;
 wire CPU_is_load_a2;
 wire CPU_is_load_a3;
 wire CPU_is_s_instr_a1;
 wire CPU_is_s_instr_a2;
 wire CPU_is_s_instr_a3;
 wire CPU_is_s_instr_a4;
 wire CPU_is_slt_a2;
 wire CPU_is_slt_a3;
 wire CPU_is_slti_a2;
 wire CPU_is_slti_a3;
 wire \CPU_pc_a2[2] ;
 wire \CPU_pc_a2[3] ;
 wire \CPU_pc_a2[4] ;
 wire \CPU_pc_a2[5] ;
 wire \CPU_rd_a2[0] ;
 wire \CPU_rd_a2[1] ;
 wire \CPU_rd_a2[2] ;
 wire \CPU_rd_a2[3] ;
 wire \CPU_rd_a2[4] ;
 wire \CPU_rd_a3[0] ;
 wire \CPU_rd_a3[1] ;
 wire \CPU_rd_a3[2] ;
 wire \CPU_rd_a3[3] ;
 wire \CPU_rd_a3[4] ;
 wire \CPU_rd_a4[0] ;
 wire \CPU_rd_a4[1] ;
 wire \CPU_rd_a4[2] ;
 wire \CPU_rd_a4[3] ;
 wire \CPU_rd_a4[4] ;
 wire \CPU_rd_a5[0] ;
 wire \CPU_rd_a5[1] ;
 wire \CPU_rd_a5[2] ;
 wire \CPU_rd_a5[3] ;
 wire \CPU_rd_a5[4] ;
 wire CPU_rd_valid_a1;
 wire CPU_rd_valid_a2;
 wire CPU_rd_valid_a3;
 wire CPU_reset_a1;
 wire CPU_reset_a2;
 wire CPU_reset_a3;
 wire CPU_reset_a4;
 wire \CPU_result_a3[2] ;
 wire \CPU_result_a3[3] ;
 wire \CPU_result_a3[4] ;
 wire \CPU_result_a3[5] ;
 wire \CPU_rf_rd_index1_a2[0] ;
 wire \CPU_rf_rd_index1_a2[1] ;
 wire \CPU_rf_rd_index1_a2[2] ;
 wire \CPU_rf_rd_index1_a2[3] ;
 wire \CPU_rf_rd_index2_a2[0] ;
 wire \CPU_rf_rd_index2_a2[1] ;
 wire \CPU_rf_rd_index2_a2[2] ;
 wire \CPU_rf_rd_index2_a2[3] ;
 wire \CPU_src1_value_a2[0] ;
 wire \CPU_src1_value_a2[10] ;
 wire \CPU_src1_value_a2[11] ;
 wire \CPU_src1_value_a2[12] ;
 wire \CPU_src1_value_a2[13] ;
 wire \CPU_src1_value_a2[14] ;
 wire \CPU_src1_value_a2[15] ;
 wire \CPU_src1_value_a2[16] ;
 wire \CPU_src1_value_a2[17] ;
 wire \CPU_src1_value_a2[18] ;
 wire \CPU_src1_value_a2[19] ;
 wire \CPU_src1_value_a2[1] ;
 wire \CPU_src1_value_a2[20] ;
 wire \CPU_src1_value_a2[21] ;
 wire \CPU_src1_value_a2[22] ;
 wire \CPU_src1_value_a2[23] ;
 wire \CPU_src1_value_a2[24] ;
 wire \CPU_src1_value_a2[25] ;
 wire \CPU_src1_value_a2[26] ;
 wire \CPU_src1_value_a2[27] ;
 wire \CPU_src1_value_a2[28] ;
 wire \CPU_src1_value_a2[29] ;
 wire \CPU_src1_value_a2[2] ;
 wire \CPU_src1_value_a2[30] ;
 wire \CPU_src1_value_a2[31] ;
 wire \CPU_src1_value_a2[3] ;
 wire \CPU_src1_value_a2[4] ;
 wire \CPU_src1_value_a2[5] ;
 wire \CPU_src1_value_a2[6] ;
 wire \CPU_src1_value_a2[7] ;
 wire \CPU_src1_value_a2[8] ;
 wire \CPU_src1_value_a2[9] ;
 wire \CPU_src1_value_a3[0] ;
 wire \CPU_src1_value_a3[10] ;
 wire \CPU_src1_value_a3[11] ;
 wire \CPU_src1_value_a3[12] ;
 wire \CPU_src1_value_a3[13] ;
 wire \CPU_src1_value_a3[14] ;
 wire \CPU_src1_value_a3[15] ;
 wire \CPU_src1_value_a3[16] ;
 wire \CPU_src1_value_a3[17] ;
 wire \CPU_src1_value_a3[18] ;
 wire \CPU_src1_value_a3[19] ;
 wire \CPU_src1_value_a3[1] ;
 wire \CPU_src1_value_a3[20] ;
 wire \CPU_src1_value_a3[21] ;
 wire \CPU_src1_value_a3[22] ;
 wire \CPU_src1_value_a3[23] ;
 wire \CPU_src1_value_a3[24] ;
 wire \CPU_src1_value_a3[25] ;
 wire \CPU_src1_value_a3[26] ;
 wire \CPU_src1_value_a3[27] ;
 wire \CPU_src1_value_a3[28] ;
 wire \CPU_src1_value_a3[29] ;
 wire \CPU_src1_value_a3[2] ;
 wire \CPU_src1_value_a3[30] ;
 wire \CPU_src1_value_a3[31] ;
 wire \CPU_src1_value_a3[3] ;
 wire \CPU_src1_value_a3[4] ;
 wire \CPU_src1_value_a3[5] ;
 wire \CPU_src1_value_a3[6] ;
 wire \CPU_src1_value_a3[7] ;
 wire \CPU_src1_value_a3[8] ;
 wire \CPU_src1_value_a3[9] ;
 wire \CPU_src2_value_a2[0] ;
 wire \CPU_src2_value_a2[10] ;
 wire \CPU_src2_value_a2[11] ;
 wire \CPU_src2_value_a2[12] ;
 wire \CPU_src2_value_a2[13] ;
 wire \CPU_src2_value_a2[14] ;
 wire \CPU_src2_value_a2[15] ;
 wire \CPU_src2_value_a2[16] ;
 wire \CPU_src2_value_a2[17] ;
 wire \CPU_src2_value_a2[18] ;
 wire \CPU_src2_value_a2[19] ;
 wire \CPU_src2_value_a2[1] ;
 wire \CPU_src2_value_a2[20] ;
 wire \CPU_src2_value_a2[21] ;
 wire \CPU_src2_value_a2[22] ;
 wire \CPU_src2_value_a2[23] ;
 wire \CPU_src2_value_a2[24] ;
 wire \CPU_src2_value_a2[25] ;
 wire \CPU_src2_value_a2[26] ;
 wire \CPU_src2_value_a2[27] ;
 wire \CPU_src2_value_a2[28] ;
 wire \CPU_src2_value_a2[29] ;
 wire \CPU_src2_value_a2[2] ;
 wire \CPU_src2_value_a2[30] ;
 wire \CPU_src2_value_a2[31] ;
 wire \CPU_src2_value_a2[3] ;
 wire \CPU_src2_value_a2[4] ;
 wire \CPU_src2_value_a2[5] ;
 wire \CPU_src2_value_a2[6] ;
 wire \CPU_src2_value_a2[7] ;
 wire \CPU_src2_value_a2[8] ;
 wire \CPU_src2_value_a2[9] ;
 wire \CPU_src2_value_a3[0] ;
 wire \CPU_src2_value_a3[10] ;
 wire \CPU_src2_value_a3[11] ;
 wire \CPU_src2_value_a3[12] ;
 wire \CPU_src2_value_a3[13] ;
 wire \CPU_src2_value_a3[14] ;
 wire \CPU_src2_value_a3[15] ;
 wire \CPU_src2_value_a3[16] ;
 wire \CPU_src2_value_a3[17] ;
 wire \CPU_src2_value_a3[18] ;
 wire \CPU_src2_value_a3[19] ;
 wire \CPU_src2_value_a3[1] ;
 wire \CPU_src2_value_a3[20] ;
 wire \CPU_src2_value_a3[21] ;
 wire \CPU_src2_value_a3[22] ;
 wire \CPU_src2_value_a3[23] ;
 wire \CPU_src2_value_a3[24] ;
 wire \CPU_src2_value_a3[25] ;
 wire \CPU_src2_value_a3[26] ;
 wire \CPU_src2_value_a3[27] ;
 wire \CPU_src2_value_a3[28] ;
 wire \CPU_src2_value_a3[29] ;
 wire \CPU_src2_value_a3[2] ;
 wire \CPU_src2_value_a3[30] ;
 wire \CPU_src2_value_a3[31] ;
 wire \CPU_src2_value_a3[3] ;
 wire \CPU_src2_value_a3[4] ;
 wire \CPU_src2_value_a3[5] ;
 wire \CPU_src2_value_a3[6] ;
 wire \CPU_src2_value_a3[7] ;
 wire \CPU_src2_value_a3[8] ;
 wire \CPU_src2_value_a3[9] ;
 wire net533;
 wire CPU_valid_a4;
 wire CPU_valid_load_a3;
 wire CPU_valid_load_a5;
 wire CPU_valid_taken_br_a3;
 wire CPU_valid_taken_br_a4;
 wire CPU_valid_taken_br_a5;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire net535;
 wire net534;
 wire net532;
 wire _01040_;
 wire _01041_;
 wire net531;
 wire _01043_;
 wire net530;
 wire net529;
 wire _01046_;
 wire net528;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire net527;
 wire _01054_;
 wire net526;
 wire net525;
 wire net524;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire net523;
 wire net522;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire net521;
 wire net520;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire net519;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire net518;
 wire net517;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire net516;
 wire net515;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire net514;
 wire net513;
 wire net512;
 wire _01126_;
 wire _01127_;
 wire net511;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire net510;
 wire _01135_;
 wire _01136_;
 wire net509;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire net508;
 wire net507;
 wire _01162_;
 wire net506;
 wire net505;
 wire net504;
 wire _01166_;
 wire net503;
 wire net502;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire net501;
 wire _01173_;
 wire _01174_;
 wire net500;
 wire net499;
 wire _01177_;
 wire _01178_;
 wire net498;
 wire _01180_;
 wire net497;
 wire net496;
 wire net495;
 wire net494;
 wire net493;
 wire _01186_;
 wire _01187_;
 wire net492;
 wire net491;
 wire _01190_;
 wire _01191_;
 wire net490;
 wire net489;
 wire _01194_;
 wire _01195_;
 wire net488;
 wire net487;
 wire _01198_;
 wire _01199_;
 wire net486;
 wire net485;
 wire _01202_;
 wire _01203_;
 wire net484;
 wire net483;
 wire _01206_;
 wire _01207_;
 wire net482;
 wire net481;
 wire _01210_;
 wire _01211_;
 wire net480;
 wire net479;
 wire _01214_;
 wire _01215_;
 wire net478;
 wire net477;
 wire _01218_;
 wire _01219_;
 wire net476;
 wire net475;
 wire net474;
 wire _01223_;
 wire net473;
 wire _01225_;
 wire net472;
 wire net471;
 wire net470;
 wire _01229_;
 wire _01230_;
 wire net469;
 wire net468;
 wire _01233_;
 wire _01234_;
 wire net467;
 wire net466;
 wire _01237_;
 wire _01238_;
 wire net465;
 wire net464;
 wire _01241_;
 wire _01242_;
 wire net463;
 wire net462;
 wire _01245_;
 wire _01246_;
 wire net461;
 wire net460;
 wire _01249_;
 wire _01250_;
 wire net459;
 wire net458;
 wire _01253_;
 wire _01254_;
 wire net457;
 wire net456;
 wire _01257_;
 wire _01258_;
 wire net455;
 wire net454;
 wire _01261_;
 wire _01262_;
 wire net453;
 wire net452;
 wire net451;
 wire _01266_;
 wire net450;
 wire _01268_;
 wire net449;
 wire net448;
 wire net447;
 wire _01272_;
 wire _01273_;
 wire net446;
 wire net445;
 wire _01276_;
 wire _01277_;
 wire net444;
 wire net443;
 wire _01280_;
 wire _01281_;
 wire net442;
 wire net441;
 wire _01284_;
 wire _01285_;
 wire net440;
 wire net439;
 wire _01288_;
 wire _01289_;
 wire net438;
 wire net437;
 wire _01292_;
 wire _01293_;
 wire net436;
 wire net435;
 wire _01296_;
 wire _01297_;
 wire net434;
 wire net433;
 wire _01300_;
 wire _01301_;
 wire net432;
 wire net431;
 wire _01304_;
 wire _01305_;
 wire net430;
 wire net429;
 wire _01308_;
 wire _01309_;
 wire net428;
 wire net427;
 wire net426;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire net425;
 wire _01317_;
 wire net424;
 wire _01319_;
 wire net423;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire net422;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire net421;
 wire _01341_;
 wire net420;
 wire _01343_;
 wire net419;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire net418;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire net417;
 wire _01367_;
 wire net416;
 wire _01369_;
 wire net415;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire net414;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire net413;
 wire _01400_;
 wire _01401_;
 wire net412;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire net411;
 wire _01419_;
 wire net410;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire net409;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire net408;
 wire _01444_;
 wire net407;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire net406;
 wire net405;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire net404;
 wire _01474_;
 wire _01475_;
 wire net403;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire net402;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire net401;
 wire _01497_;
 wire net400;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire net399;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire net398;
 wire _01520_;
 wire net397;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire net396;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire net395;
 wire _01551_;
 wire net394;
 wire _01553_;
 wire _01554_;
 wire net393;
 wire _01556_;
 wire _01557_;
 wire net392;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire net391;
 wire _01575_;
 wire net390;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire net389;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire net388;
 wire _01598_;
 wire net387;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire net386;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire net385;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire net384;
 wire _01634_;
 wire net383;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire net382;
 wire _01649_;
 wire net381;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire net380;
 wire net379;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire net378;
 wire _01675_;
 wire net377;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire net376;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire net375;
 wire _01708_;
 wire _01709_;
 wire net374;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire net373;
 wire net372;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire net371;
 wire _01727_;
 wire net370;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire net369;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire net368;
 wire _01752_;
 wire net367;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire net366;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire net365;
 wire _01785_;
 wire _01786_;
 wire net364;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire net363;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire net362;
 wire _01809_;
 wire net361;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire net360;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire net359;
 wire _01832_;
 wire net358;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire net357;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire net356;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire net355;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire net354;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire net353;
 wire _01883_;
 wire net352;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire net351;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire net350;
 wire _01908_;
 wire net349;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire net348;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire net347;
 wire _01936_;
 wire net346;
 wire _01938_;
 wire _01939_;
 wire net345;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire net344;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire net343;
 wire _01960_;
 wire net342;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire net341;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire net340;
 wire net339;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire net338;
 wire _01987_;
 wire net337;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire net336;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire net335;
 wire _02015_;
 wire net334;
 wire _02017_;
 wire _02018_;
 wire net333;
 wire _02020_;
 wire net332;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire net331;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire net330;
 wire _02041_;
 wire net329;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire net328;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire net327;
 wire _02064_;
 wire net326;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire net325;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire net324;
 wire _02094_;
 wire net323;
 wire _02096_;
 wire _02097_;
 wire net322;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire net321;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire net320;
 wire _02118_;
 wire net319;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire net318;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire net317;
 wire _02141_;
 wire net316;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire net315;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire net314;
 wire _02171_;
 wire _02172_;
 wire net313;
 wire _02174_;
 wire net312;
 wire _02176_;
 wire net311;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire net310;
 wire _02193_;
 wire net309;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire net308;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire net307;
 wire _02218_;
 wire net306;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire net305;
 wire net304;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire net303;
 wire _02249_;
 wire net302;
 wire _02251_;
 wire _02252_;
 wire net301;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire net300;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire net299;
 wire _02271_;
 wire net298;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire net297;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire net296;
 wire _02296_;
 wire net295;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire net294;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire net293;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire net292;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire net291;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire net290;
 wire _02349_;
 wire net289;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire net288;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire net287;
 wire _02372_;
 wire net286;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire net285;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire net284;
 wire _02403_;
 wire _02404_;
 wire net283;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire net282;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire net281;
 wire _02425_;
 wire net280;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire net279;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire net278;
 wire _02448_;
 wire net277;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire net276;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire net275;
 wire net274;
 wire net273;
 wire net272;
 wire net271;
 wire net270;
 wire _02482_;
 wire _02483_;
 wire net269;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire net268;
 wire net267;
 wire _02493_;
 wire net266;
 wire net265;
 wire net264;
 wire _02497_;
 wire net263;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire net262;
 wire net261;
 wire net260;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire net259;
 wire net258;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire net257;
 wire _02562_;
 wire net256;
 wire _02564_;
 wire net255;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire net254;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire net253;
 wire net252;
 wire net251;
 wire _02586_;
 wire net250;
 wire _02588_;
 wire net249;
 wire net248;
 wire net247;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire net246;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire net245;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire net244;
 wire net243;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire net242;
 wire _02639_;
 wire net241;
 wire _02641_;
 wire net240;
 wire net239;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire net238;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire net237;
 wire net236;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire net235;
 wire net234;
 wire net233;
 wire net232;
 wire net231;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire net230;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire net229;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire net228;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire net227;
 wire _02811_;
 wire net226;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire net225;
 wire _02834_;
 wire net224;
 wire net223;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire net222;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire net221;
 wire _02884_;
 wire net220;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire net219;
 wire _02891_;
 wire net218;
 wire net217;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire net216;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire net215;
 wire _02936_;
 wire net214;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire net213;
 wire _02961_;
 wire net212;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire net211;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire net210;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire net209;
 wire net208;
 wire net207;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire net206;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire net205;
 wire _03076_;
 wire net204;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire net203;
 wire _03100_;
 wire net202;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire net201;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire net200;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire net199;
 wire net198;
 wire _03138_;
 wire _03139_;
 wire net197;
 wire net196;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire net195;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire net194;
 wire _03163_;
 wire net193;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire net192;
 wire _03191_;
 wire net191;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire net190;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire net189;
 wire _03238_;
 wire net188;
 wire net187;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire net186;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire net185;
 wire _03261_;
 wire net184;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire _03275_;
 wire net179;
 wire _03277_;
 wire _03278_;
 wire net178;
 wire _03280_;
 wire _03281_;
 wire net177;
 wire _03283_;
 wire net176;
 wire _03285_;
 wire net175;
 wire net174;
 wire net173;
 wire _03289_;
 wire net172;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire net171;
 wire _03297_;
 wire net170;
 wire _03299_;
 wire net169;
 wire net168;
 wire _03302_;
 wire net167;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire net166;
 wire _03308_;
 wire net165;
 wire _03310_;
 wire net164;
 wire _03312_;
 wire _03313_;
 wire net163;
 wire _03315_;
 wire net162;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire net161;
 wire _03321_;
 wire _03322_;
 wire net160;
 wire _03324_;
 wire _03325_;
 wire net159;
 wire _03327_;
 wire net158;
 wire _03329_;
 wire _03330_;
 wire net157;
 wire net156;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire net155;
 wire net154;
 wire _03339_;
 wire _03340_;
 wire net153;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire net152;
 wire _03346_;
 wire _03347_;
 wire net151;
 wire _03349_;
 wire _03350_;
 wire net150;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire net149;
 wire net148;
 wire net147;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire net146;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire net145;
 wire _03375_;
 wire net144;
 wire _03377_;
 wire _03378_;
 wire net143;
 wire net142;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire net141;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire net140;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire net139;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire net138;
 wire net137;
 wire net136;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire net135;
 wire _03441_;
 wire _03442_;
 wire net134;
 wire _03444_;
 wire _03445_;
 wire net133;
 wire net132;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire net131;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire net130;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire net129;
 wire net128;
 wire net127;
 wire _03500_;
 wire net126;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire net125;
 wire _03506_;
 wire net124;
 wire _03508_;
 wire _03509_;
 wire net123;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire net122;
 wire net121;
 wire _03519_;
 wire net120;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire net119;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire net118;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire net117;
 wire net116;
 wire net115;
 wire _03563_;
 wire _03564_;
 wire net114;
 wire _03566_;
 wire _03567_;
 wire clknet_4_15_0_clk;
 wire _03569_;
 wire _03570_;
 wire clknet_4_14_0_clk;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire clknet_4_13_0_clk;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire clknet_4_12_0_clk;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire clknet_4_11_0_clk;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire clknet_4_10_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_8_0_clk;
 wire _03626_;
 wire _03627_;
 wire clknet_4_7_0_clk;
 wire _03629_;
 wire _03630_;
 wire clknet_4_6_0_clk;
 wire _03632_;
 wire _03633_;
 wire clknet_4_5_0_clk;
 wire clknet_4_4_0_clk;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire clknet_4_3_0_clk;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire clknet_4_2_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_0_0_clk;
 wire _03689_;
 wire clknet_0_clk;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire clknet_leaf_122_clk;
 wire _03695_;
 wire clknet_leaf_121_clk;
 wire _03697_;
 wire _03698_;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_118_clk;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire clknet_leaf_117_clk;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire clknet_leaf_116_clk;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire clknet_leaf_115_clk;
 wire _03749_;
 wire _03750_;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_112_clk;
 wire _03754_;
 wire _03755_;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_110_clk;
 wire _03758_;
 wire _03759_;
 wire clknet_leaf_109_clk;
 wire _03761_;
 wire _03762_;
 wire clknet_leaf_108_clk;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire clknet_leaf_107_clk;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire clknet_leaf_106_clk;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire clknet_leaf_105_clk;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_102_clk;
 wire _03821_;
 wire _03822_;
 wire clknet_leaf_101_clk;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire clknet_leaf_100_clk;
 wire _03828_;
 wire clknet_leaf_99_clk;
 wire _03830_;
 wire _03831_;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_96_clk;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire clknet_leaf_95_clk;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire clknet_leaf_94_clk;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_91_clk;
 wire _03886_;
 wire _03887_;
 wire clknet_leaf_90_clk;
 wire _03889_;
 wire _03890_;
 wire clknet_leaf_89_clk;
 wire _03892_;
 wire _03893_;
 wire clknet_leaf_88_clk;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire clknet_leaf_87_clk;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_83_clk;
 wire _03948_;
 wire clknet_leaf_82_clk;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire clknet_leaf_81_clk;
 wire _03954_;
 wire clknet_leaf_80_clk;
 wire _03956_;
 wire _03957_;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_76_clk;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_73_clk;
 wire _04010_;
 wire _04011_;
 wire clknet_leaf_72_clk;
 wire _04013_;
 wire clknet_leaf_71_clk;
 wire _04015_;
 wire clknet_leaf_70_clk;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire clknet_leaf_69_clk;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire clknet_leaf_68_clk;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire clknet_leaf_67_clk;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_64_clk;
 wire _04072_;
 wire clknet_leaf_63_clk;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire clknet_leaf_62_clk;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_58_clk;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire clknet_leaf_57_clk;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_54_clk;
 wire _04135_;
 wire _04136_;
 wire clknet_leaf_53_clk;
 wire _04138_;
 wire _04139_;
 wire clknet_leaf_52_clk;
 wire _04141_;
 wire _04142_;
 wire clknet_leaf_51_clk;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_49_clk;
 wire _04227_;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_47_clk;
 wire _04230_;
 wire _04231_;
 wire clknet_leaf_46_clk;
 wire _04233_;
 wire _04234_;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_44_clk;
 wire _04237_;
 wire clknet_leaf_43_clk;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_41_clk;
 wire _04244_;
 wire _04245_;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_39_clk;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire clknet_leaf_38_clk;
 wire _04252_;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_36_clk;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire clknet_leaf_35_clk;
 wire _04260_;
 wire clknet_leaf_34_clk;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire clknet_leaf_33_clk;
 wire _04266_;
 wire clknet_leaf_32_clk;
 wire _04268_;
 wire _04269_;
 wire clknet_leaf_31_clk;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire clknet_leaf_30_clk;
 wire _04275_;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_28_clk;
 wire _04278_;
 wire _04279_;
 wire clknet_leaf_27_clk;
 wire _04281_;
 wire clknet_leaf_26_clk;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_22_clk;
 wire _04297_;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire _04300_;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire _04303_;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire _04306_;
 wire _04307_;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire _04310_;
 wire _04311_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire _04314_;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_9_clk;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire clknet_leaf_8_clk;
 wire _04322_;
 wire clknet_leaf_7_clk;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire _04333_;
 wire clknet_leaf_4_clk;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire clknet_leaf_3_clk;
 wire _04341_;
 wire clknet_leaf_2_clk;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire clknet_leaf_1_clk;
 wire _04350_;
 wire net113;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire net112;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire net111;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire net110;
 wire _04377_;
 wire net109;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire net108;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire net107;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire net106;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire net105;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire _04692_;
 wire net100;
 wire net99;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire net98;
 wire net97;
 wire _04700_;
 wire net96;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire net95;
 wire _04707_;
 wire net94;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire net93;
 wire _04713_;
 wire net92;
 wire _04715_;
 wire _04716_;
 wire net91;
 wire _04718_;
 wire _04719_;
 wire net90;
 wire net89;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire net88;
 wire _04726_;
 wire net87;
 wire net86;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire net85;
 wire net84;
 wire _04736_;
 wire net83;
 wire net82;
 wire _04739_;
 wire _04740_;
 wire net81;
 wire _04742_;
 wire net80;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire _04757_;
 wire net75;
 wire net74;
 wire _04760_;
 wire net73;
 wire net72;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire net71;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire net70;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire net69;
 wire _04775_;
 wire net68;
 wire _04777_;
 wire net67;
 wire _04779_;
 wire net66;
 wire _04781_;
 wire net65;
 wire _04783_;
 wire _04784_;
 wire net64;
 wire net63;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire net62;
 wire net61;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire net60;
 wire net59;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire net58;
 wire net57;
 wire _04807_;
 wire net56;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire net55;
 wire _04817_;
 wire _04818_;
 wire net54;
 wire net53;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire net52;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire net51;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire net50;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire net49;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire net48;
 wire _04858_;
 wire _04859_;
 wire net47;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire net46;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire net45;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire net44;
 wire net43;
 wire net42;
 wire _05146_;
 wire net41;
 wire net40;
 wire _05149_;
 wire net39;
 wire net38;
 wire _05152_;
 wire net37;
 wire net36;
 wire _05155_;
 wire _05156_;
 wire net35;
 wire net34;
 wire _05159_;
 wire net33;
 wire net32;
 wire _05162_;
 wire net31;
 wire net30;
 wire net29;
 wire _05166_;
 wire net28;
 wire net27;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire net26;
 wire _05173_;
 wire net25;
 wire net24;
 wire _05176_;
 wire net23;
 wire net22;
 wire _05179_;
 wire _05180_;
 wire net21;
 wire _05182_;
 wire _05183_;
 wire net20;
 wire _05185_;
 wire net19;
 wire _05187_;
 wire _05188_;
 wire net18;
 wire _05190_;
 wire _05191_;
 wire net17;
 wire _05193_;
 wire net16;
 wire net15;
 wire _05196_;
 wire _05197_;
 wire net14;
 wire _05199_;
 wire _05200_;
 wire net13;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire net12;
 wire _05207_;
 wire net11;
 wire net10;
 wire _05210_;
 wire net9;
 wire net8;
 wire _05213_;
 wire _05214_;
 wire net7;
 wire _05216_;
 wire _05217_;
 wire net6;
 wire _05219_;
 wire net5;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire net4;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire net3;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire net2;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire net1;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire clknet_leaf_0_clk;
 wire \w_CPU_dmem_rd_data_a4[0] ;
 wire \w_CPU_dmem_rd_data_a4[10] ;
 wire \w_CPU_dmem_rd_data_a4[11] ;
 wire \w_CPU_dmem_rd_data_a4[12] ;
 wire \w_CPU_dmem_rd_data_a4[13] ;
 wire \w_CPU_dmem_rd_data_a4[14] ;
 wire \w_CPU_dmem_rd_data_a4[15] ;
 wire \w_CPU_dmem_rd_data_a4[16] ;
 wire \w_CPU_dmem_rd_data_a4[17] ;
 wire \w_CPU_dmem_rd_data_a4[18] ;
 wire \w_CPU_dmem_rd_data_a4[19] ;
 wire \w_CPU_dmem_rd_data_a4[1] ;
 wire \w_CPU_dmem_rd_data_a4[20] ;
 wire \w_CPU_dmem_rd_data_a4[21] ;
 wire \w_CPU_dmem_rd_data_a4[22] ;
 wire \w_CPU_dmem_rd_data_a4[23] ;
 wire \w_CPU_dmem_rd_data_a4[24] ;
 wire \w_CPU_dmem_rd_data_a4[25] ;
 wire \w_CPU_dmem_rd_data_a4[26] ;
 wire \w_CPU_dmem_rd_data_a4[27] ;
 wire \w_CPU_dmem_rd_data_a4[28] ;
 wire \w_CPU_dmem_rd_data_a4[29] ;
 wire \w_CPU_dmem_rd_data_a4[2] ;
 wire \w_CPU_dmem_rd_data_a4[30] ;
 wire \w_CPU_dmem_rd_data_a4[31] ;
 wire \w_CPU_dmem_rd_data_a4[3] ;
 wire \w_CPU_dmem_rd_data_a4[4] ;
 wire \w_CPU_dmem_rd_data_a4[5] ;
 wire \w_CPU_dmem_rd_data_a4[6] ;
 wire \w_CPU_dmem_rd_data_a4[7] ;
 wire \w_CPU_dmem_rd_data_a4[8] ;
 wire \w_CPU_dmem_rd_data_a4[9] ;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;

 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][0]$_SDFFE_PP0P_  (.D(net849),
    .Q(\CPU_Dmem_value_a5[0][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][10]$_SDFFE_PP0P_  (.D(net501),
    .Q(\CPU_Dmem_value_a5[0][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][11]$_SDFFE_PP0P_  (.D(net300),
    .Q(\CPU_Dmem_value_a5[0][11] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][12]$_SDFFE_PP0P_  (.D(net372),
    .Q(\CPU_Dmem_value_a5[0][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][13]$_SDFFE_PP0P_  (.D(net538),
    .Q(\CPU_Dmem_value_a5[0][13] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][14]$_SDFFE_PP0P_  (.D(net316),
    .Q(\CPU_Dmem_value_a5[0][14] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][15]$_SDFFE_PP0P_  (.D(net473),
    .Q(\CPU_Dmem_value_a5[0][15] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][16]$_SDFFE_PP0P_  (.D(net1163),
    .Q(\CPU_Dmem_value_a5[0][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][17]$_SDFFE_PP0P_  (.D(net742),
    .Q(\CPU_Dmem_value_a5[0][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][18]$_SDFFE_PP0P_  (.D(net1019),
    .Q(\CPU_Dmem_value_a5[0][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][19]$_SDFFE_PP0P_  (.D(net544),
    .Q(\CPU_Dmem_value_a5[0][19] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][1]$_SDFFE_PP0P_  (.D(net388),
    .Q(\CPU_Dmem_value_a5[0][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][20]$_SDFFE_PP0P_  (.D(net647),
    .Q(\CPU_Dmem_value_a5[0][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][21]$_SDFFE_PP0P_  (.D(net839),
    .Q(\CPU_Dmem_value_a5[0][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][22]$_SDFFE_PP0P_  (.D(net1078),
    .Q(\CPU_Dmem_value_a5[0][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][23]$_SDFFE_PP0P_  (.D(net776),
    .Q(\CPU_Dmem_value_a5[0][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][24]$_SDFFE_PP0P_  (.D(net384),
    .Q(\CPU_Dmem_value_a5[0][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][25]$_SDFFE_PP0P_  (.D(net554),
    .Q(\CPU_Dmem_value_a5[0][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][26]$_SDFFE_PP0P_  (.D(net1076),
    .Q(\CPU_Dmem_value_a5[0][26] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][27]$_SDFFE_PP0P_  (.D(net845),
    .Q(\CPU_Dmem_value_a5[0][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][28]$_SDFFE_PP0P_  (.D(net754),
    .Q(\CPU_Dmem_value_a5[0][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][29]$_SDFFE_PP0P_  (.D(net370),
    .Q(\CPU_Dmem_value_a5[0][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][2]$_SDFFE_PP0P_  (.D(net400),
    .Q(\CPU_Dmem_value_a5[0][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][30]$_SDFFE_PP0P_  (.D(net1084),
    .Q(\CPU_Dmem_value_a5[0][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][31]$_SDFFE_PP0P_  (.D(net451),
    .Q(\CPU_Dmem_value_a5[0][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][3]$_SDFFE_PP0P_  (.D(net993),
    .Q(\CPU_Dmem_value_a5[0][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][4]$_SDFFE_PP0P_  (.D(net730),
    .Q(\CPU_Dmem_value_a5[0][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][5]$_SDFFE_PP0P_  (.D(net489),
    .Q(\CPU_Dmem_value_a5[0][5] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][6]$_SDFFE_PP0P_  (.D(net891),
    .Q(\CPU_Dmem_value_a5[0][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][7]$_SDFFE_PP0P_  (.D(net790),
    .Q(\CPU_Dmem_value_a5[0][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][8]$_SDFFE_PP0P_  (.D(net540),
    .Q(\CPU_Dmem_value_a5[0][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[0][9]$_SDFFE_PP0P_  (.D(net1382),
    .Q(\CPU_Dmem_value_a5[0][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][0]$_SDFFE_PP0P_  (.D(net786),
    .Q(\CPU_Dmem_value_a5[10][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][10]$_SDFFE_PP0P_  (.D(net457),
    .Q(\CPU_Dmem_value_a5[10][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][11]$_SDFFE_PP0P_  (.D(net534),
    .Q(\CPU_Dmem_value_a5[10][11] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][12]$_SDFFE_PP0P_  (.D(net242),
    .Q(\CPU_Dmem_value_a5[10][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][13]$_SDFFE_PP0P_  (.D(net910),
    .Q(\CPU_Dmem_value_a5[10][13] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][14]$_SDFFE_PP0P_  (.D(net230),
    .Q(\CPU_Dmem_value_a5[10][14] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][15]$_SDFFE_PP0P_  (.D(net953),
    .Q(\CPU_Dmem_value_a5[10][15] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][16]$_SDFFE_PP0P_  (.D(net943),
    .Q(\CPU_Dmem_value_a5[10][16] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][17]$_SDFFE_PP0P_  (.D(net447),
    .Q(\CPU_Dmem_value_a5[10][17] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][18]$_SDFFE_PP0P_  (.D(net344),
    .Q(\CPU_Dmem_value_a5[10][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][19]$_SDFFE_PP0P_  (.D(net1207),
    .Q(\CPU_Dmem_value_a5[10][19] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][1]$_SDFFE_PP1P_  (.D(net1074),
    .Q(\CPU_Dmem_value_a5[10][1] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][20]$_SDFFE_PP0P_  (.D(net479),
    .Q(\CPU_Dmem_value_a5[10][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][21]$_SDFFE_PP0P_  (.D(net350),
    .Q(\CPU_Dmem_value_a5[10][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][22]$_SDFFE_PP0P_  (.D(net1102),
    .Q(\CPU_Dmem_value_a5[10][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][23]$_SDFFE_PP0P_  (.D(net820),
    .Q(\CPU_Dmem_value_a5[10][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][24]$_SDFFE_PP0P_  (.D(net556),
    .Q(\CPU_Dmem_value_a5[10][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][25]$_SDFFE_PP0P_  (.D(net481),
    .Q(\CPU_Dmem_value_a5[10][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][26]$_SDFFE_PP0P_  (.D(net947),
    .Q(\CPU_Dmem_value_a5[10][26] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][27]$_SDFFE_PP0P_  (.D(net851),
    .Q(\CPU_Dmem_value_a5[10][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][28]$_SDFFE_PP0P_  (.D(net985),
    .Q(\CPU_Dmem_value_a5[10][28] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][29]$_SDFFE_PP0P_  (.D(net586),
    .Q(\CPU_Dmem_value_a5[10][29] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][2]$_SDFFE_PP0P_  (.D(net467),
    .Q(\CPU_Dmem_value_a5[10][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][30]$_SDFFE_PP0P_  (.D(net483),
    .Q(\CPU_Dmem_value_a5[10][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][31]$_SDFFE_PP0P_  (.D(net904),
    .Q(\CPU_Dmem_value_a5[10][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][3]$_SDFFE_PP1P_  (.D(net1128),
    .Q(\CPU_Dmem_value_a5[10][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][4]$_SDFFE_PP0P_  (.D(net921),
    .Q(\CPU_Dmem_value_a5[10][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][5]$_SDFFE_PP0P_  (.D(net362),
    .Q(\CPU_Dmem_value_a5[10][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][6]$_SDFFE_PP0P_  (.D(net951),
    .Q(\CPU_Dmem_value_a5[10][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][7]$_SDFFE_PP0P_  (.D(net1035),
    .Q(\CPU_Dmem_value_a5[10][7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][8]$_SDFFE_PP0P_  (.D(net493),
    .Q(\CPU_Dmem_value_a5[10][8] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[10][9]$_SDFFE_PP0P_  (.D(net455),
    .Q(\CPU_Dmem_value_a5[10][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][0]$_SDFFE_PP1P_  (.D(net981),
    .Q(\CPU_Dmem_value_a5[11][0] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][10]$_SDFFE_PP0P_  (.D(net394),
    .Q(\CPU_Dmem_value_a5[11][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][11]$_SDFFE_PP0P_  (.D(net615),
    .Q(\CPU_Dmem_value_a5[11][11] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][12]$_SDFFE_PP0P_  (.D(net356),
    .Q(\CPU_Dmem_value_a5[11][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][13]$_SDFFE_PP0P_  (.D(net348),
    .Q(\CPU_Dmem_value_a5[11][13] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][14]$_SDFFE_PP0P_  (.D(net867),
    .Q(\CPU_Dmem_value_a5[11][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][15]$_SDFFE_PP0P_  (.D(net633),
    .Q(\CPU_Dmem_value_a5[11][15] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][16]$_SDFFE_PP0P_  (.D(net979),
    .Q(\CPU_Dmem_value_a5[11][16] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][17]$_SDFFE_PP0P_  (.D(net530),
    .Q(\CPU_Dmem_value_a5[11][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][18]$_SDFFE_PP0P_  (.D(net603),
    .Q(\CPU_Dmem_value_a5[11][18] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][19]$_SDFFE_PP0P_  (.D(net412),
    .Q(\CPU_Dmem_value_a5[11][19] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][1]$_SDFFE_PP1P_  (.D(net1209),
    .Q(\CPU_Dmem_value_a5[11][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][20]$_SDFFE_PP0P_  (.D(net336),
    .Q(\CPU_Dmem_value_a5[11][20] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][21]$_SDFFE_PP0P_  (.D(net681),
    .Q(\CPU_Dmem_value_a5[11][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][22]$_SDFFE_PP0P_  (.D(net1023),
    .Q(\CPU_Dmem_value_a5[11][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][23]$_SDFFE_PP0P_  (.D(net885),
    .Q(\CPU_Dmem_value_a5[11][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][24]$_SDFFE_PP0P_  (.D(net1009),
    .Q(\CPU_Dmem_value_a5[11][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][25]$_SDFFE_PP0P_  (.D(net1058),
    .Q(\CPU_Dmem_value_a5[11][25] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][26]$_SDFFE_PP0P_  (.D(net941),
    .Q(\CPU_Dmem_value_a5[11][26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][27]$_SDFFE_PP0P_  (.D(net897),
    .Q(\CPU_Dmem_value_a5[11][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][28]$_SDFFE_PP0P_  (.D(net443),
    .Q(\CPU_Dmem_value_a5[11][28] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][29]$_SDFFE_PP0P_  (.D(net560),
    .Q(\CPU_Dmem_value_a5[11][29] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][2]$_SDFFE_PP0P_  (.D(net806),
    .Q(\CPU_Dmem_value_a5[11][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][30]$_SDFFE_PP0P_  (.D(net408),
    .Q(\CPU_Dmem_value_a5[11][30] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][31]$_SDFFE_PP0P_  (.D(net621),
    .Q(\CPU_Dmem_value_a5[11][31] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][3]$_SDFFE_PP1P_  (.D(net1060),
    .Q(\CPU_Dmem_value_a5[11][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][4]$_SDFFE_PP0P_  (.D(net746),
    .Q(\CPU_Dmem_value_a5[11][4] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][5]$_SDFFE_PP0P_  (.D(net1175),
    .Q(\CPU_Dmem_value_a5[11][5] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][6]$_SDFFE_PP0P_  (.D(net631),
    .Q(\CPU_Dmem_value_a5[11][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][7]$_SDFFE_PP0P_  (.D(net969),
    .Q(\CPU_Dmem_value_a5[11][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][8]$_SDFFE_PP0P_  (.D(net673),
    .Q(\CPU_Dmem_value_a5[11][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[11][9]$_SDFFE_PP0P_  (.D(net1330),
    .Q(\CPU_Dmem_value_a5[11][9] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][0]$_SDFFE_PP0P_  (.D(net552),
    .Q(\CPU_Dmem_value_a5[12][0] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][10]$_SDFFE_PP0P_  (.D(net438),
    .Q(\CPU_Dmem_value_a5[12][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][11]$_SDFFE_PP0P_  (.D(net835),
    .Q(\CPU_Dmem_value_a5[12][11] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][12]$_SDFFE_PP0P_  (.D(net1106),
    .Q(\CPU_Dmem_value_a5[12][12] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][13]$_SDFFE_PP0P_  (.D(net330),
    .Q(\CPU_Dmem_value_a5[12][13] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][14]$_SDFFE_PP0P_  (.D(net558),
    .Q(\CPU_Dmem_value_a5[12][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][15]$_SDFFE_PP0P_  (.D(net1122),
    .Q(\CPU_Dmem_value_a5[12][15] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][16]$_SDFFE_PP0P_  (.D(net802),
    .Q(\CPU_Dmem_value_a5[12][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][17]$_SDFFE_PP0P_  (.D(net461),
    .Q(\CPU_Dmem_value_a5[12][17] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][18]$_SDFFE_PP0P_  (.D(net701),
    .Q(\CPU_Dmem_value_a5[12][18] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][19]$_SDFFE_PP0P_  (.D(net410),
    .Q(\CPU_Dmem_value_a5[12][19] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][1]$_SDFFE_PP0P_  (.D(net788),
    .Q(\CPU_Dmem_value_a5[12][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][20]$_SDFFE_PP0P_  (.D(net625),
    .Q(\CPU_Dmem_value_a5[12][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][21]$_SDFFE_PP0P_  (.D(net477),
    .Q(\CPU_Dmem_value_a5[12][21] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][22]$_SDFFE_PP0P_  (.D(net857),
    .Q(\CPU_Dmem_value_a5[12][22] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][23]$_SDFFE_PP0P_  (.D(net923),
    .Q(\CPU_Dmem_value_a5[12][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][24]$_SDFFE_PP0P_  (.D(net1110),
    .Q(\CPU_Dmem_value_a5[12][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][25]$_SDFFE_PP0P_  (.D(net254),
    .Q(\CPU_Dmem_value_a5[12][25] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][26]$_SDFFE_PP0P_  (.D(net881),
    .Q(\CPU_Dmem_value_a5[12][26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][27]$_SDFFE_PP0P_  (.D(net453),
    .Q(\CPU_Dmem_value_a5[12][27] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][28]$_SDFFE_PP0P_  (.D(net824),
    .Q(\CPU_Dmem_value_a5[12][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][29]$_SDFFE_PP0P_  (.D(net780),
    .Q(\CPU_Dmem_value_a5[12][29] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][2]$_SDFFE_PP1P_  (.D(net1220),
    .Q(\CPU_Dmem_value_a5[12][2] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][30]$_SDFFE_PP0P_  (.D(net683),
    .Q(\CPU_Dmem_value_a5[12][30] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][31]$_SDFFE_PP0P_  (.D(net1534),
    .Q(\CPU_Dmem_value_a5[12][31] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][3]$_SDFFE_PP1P_  (.D(net1232),
    .Q(\CPU_Dmem_value_a5[12][3] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][4]$_SDFFE_PP0P_  (.D(net518),
    .Q(\CPU_Dmem_value_a5[12][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][5]$_SDFFE_PP0P_  (.D(net1345),
    .Q(\CPU_Dmem_value_a5[12][5] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][6]$_SDFFE_PP0P_  (.D(net1203),
    .Q(\CPU_Dmem_value_a5[12][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][7]$_SDFFE_PP0P_  (.D(net629),
    .Q(\CPU_Dmem_value_a5[12][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][8]$_SDFFE_PP0P_  (.D(net762),
    .Q(\CPU_Dmem_value_a5[12][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[12][9]$_SDFFE_PP0P_  (.D(net1194),
    .Q(\CPU_Dmem_value_a5[12][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][0]$_SDFFE_PP1P_  (.D(net1252),
    .Q(\CPU_Dmem_value_a5[13][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][10]$_SDFFE_PP0P_  (.D(net1130),
    .Q(\CPU_Dmem_value_a5[13][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][11]$_SDFFE_PP0P_  (.D(net671),
    .Q(\CPU_Dmem_value_a5[13][11] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][12]$_SDFFE_PP0P_  (.D(net459),
    .Q(\CPU_Dmem_value_a5[13][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][13]$_SDFFE_PP0P_  (.D(net1112),
    .Q(\CPU_Dmem_value_a5[13][13] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][14]$_SDFFE_PP0P_  (.D(net250),
    .Q(\CPU_Dmem_value_a5[13][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][15]$_SDFFE_PP0P_  (.D(net695),
    .Q(\CPU_Dmem_value_a5[13][15] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][16]$_SDFFE_PP0P_  (.D(net712),
    .Q(\CPU_Dmem_value_a5[13][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][17]$_SDFFE_PP0P_  (.D(net657),
    .Q(\CPU_Dmem_value_a5[13][17] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][18]$_SDFFE_PP0P_  (.D(net738),
    .Q(\CPU_Dmem_value_a5[13][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][19]$_SDFFE_PP0P_  (.D(net342),
    .Q(\CPU_Dmem_value_a5[13][19] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][1]$_SDFFE_PP0P_  (.D(net506),
    .Q(\CPU_Dmem_value_a5[13][1] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][20]$_SDFFE_PP0P_  (.D(net1148),
    .Q(\CPU_Dmem_value_a5[13][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][21]$_SDFFE_PP0P_  (.D(net877),
    .Q(\CPU_Dmem_value_a5[13][21] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][22]$_SDFFE_PP0P_  (.D(net810),
    .Q(\CPU_Dmem_value_a5[13][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][23]$_SDFFE_PP0P_  (.D(net902),
    .Q(\CPU_Dmem_value_a5[13][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][24]$_SDFFE_PP0P_  (.D(net1094),
    .Q(\CPU_Dmem_value_a5[13][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][25]$_SDFFE_PP0P_  (.D(net366),
    .Q(\CPU_Dmem_value_a5[13][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][26]$_SDFFE_PP0P_  (.D(net432),
    .Q(\CPU_Dmem_value_a5[13][26] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][27]$_SDFFE_PP0P_  (.D(net816),
    .Q(\CPU_Dmem_value_a5[13][27] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][28]$_SDFFE_PP0P_  (.D(net1015),
    .Q(\CPU_Dmem_value_a5[13][28] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][29]$_SDFFE_PP0P_  (.D(net814),
    .Q(\CPU_Dmem_value_a5[13][29] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][2]$_SDFFE_PP1P_  (.D(net1349),
    .Q(\CPU_Dmem_value_a5[13][2] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][30]$_SDFFE_PP0P_  (.D(net1047),
    .Q(\CPU_Dmem_value_a5[13][30] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][31]$_SDFFE_PP0P_  (.D(net914),
    .Q(\CPU_Dmem_value_a5[13][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][3]$_SDFFE_PP1P_  (.D(net1265),
    .Q(\CPU_Dmem_value_a5[13][3] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][4]$_SDFFE_PP0P_  (.D(net655),
    .Q(\CPU_Dmem_value_a5[13][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][5]$_SDFFE_PP0P_  (.D(net995),
    .Q(\CPU_Dmem_value_a5[13][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][6]$_SDFFE_PP0P_  (.D(net292),
    .Q(\CPU_Dmem_value_a5[13][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][7]$_SDFFE_PP0P_  (.D(net679),
    .Q(\CPU_Dmem_value_a5[13][7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][8]$_SDFFE_PP0P_  (.D(net1153),
    .Q(\CPU_Dmem_value_a5[13][8] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[13][9]$_SDFFE_PP0P_  (.D(net1247),
    .Q(\CPU_Dmem_value_a5[13][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][0]$_SDFFE_PP0P_  (.D(net520),
    .Q(\CPU_Dmem_value_a5[14][0] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][10]$_SDFFE_PP0P_  (.D(net352),
    .Q(\CPU_Dmem_value_a5[14][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][11]$_SDFFE_PP0P_  (.D(net784),
    .Q(\CPU_Dmem_value_a5[14][11] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][12]$_SDFFE_PP0P_  (.D(net778),
    .Q(\CPU_Dmem_value_a5[14][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][13]$_SDFFE_PP0P_  (.D(net607),
    .Q(\CPU_Dmem_value_a5[14][13] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][14]$_SDFFE_PP0P_  (.D(net965),
    .Q(\CPU_Dmem_value_a5[14][14] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][15]$_SDFFE_PP0P_  (.D(net516),
    .Q(\CPU_Dmem_value_a5[14][15] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][16]$_SDFFE_PP0P_  (.D(net1088),
    .Q(\CPU_Dmem_value_a5[14][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][17]$_SDFFE_PP0P_  (.D(net276),
    .Q(\CPU_Dmem_value_a5[14][17] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][18]$_SDFFE_PP0P_  (.D(net697),
    .Q(\CPU_Dmem_value_a5[14][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][19]$_SDFFE_PP0P_  (.D(net358),
    .Q(\CPU_Dmem_value_a5[14][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][1]$_SDFFE_PP1P_  (.D(net1301),
    .Q(\CPU_Dmem_value_a5[14][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][20]$_SDFFE_PP0P_  (.D(net1062),
    .Q(\CPU_Dmem_value_a5[14][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][21]$_SDFFE_PP0P_  (.D(net576),
    .Q(\CPU_Dmem_value_a5[14][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][22]$_SDFFE_PP0P_  (.D(net228),
    .Q(\CPU_Dmem_value_a5[14][22] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][23]$_SDFFE_PP0P_  (.D(net665),
    .Q(\CPU_Dmem_value_a5[14][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][24]$_SDFFE_PP0P_  (.D(net782),
    .Q(\CPU_Dmem_value_a5[14][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][25]$_SDFFE_PP0P_  (.D(net1013),
    .Q(\CPU_Dmem_value_a5[14][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][26]$_SDFFE_PP0P_  (.D(net258),
    .Q(\CPU_Dmem_value_a5[14][26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][27]$_SDFFE_PP0P_  (.D(net590),
    .Q(\CPU_Dmem_value_a5[14][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][28]$_SDFFE_PP0P_  (.D(net714),
    .Q(\CPU_Dmem_value_a5[14][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][29]$_SDFFE_PP0P_  (.D(net542),
    .Q(\CPU_Dmem_value_a5[14][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][2]$_SDFFE_PP1P_  (.D(net1222),
    .Q(\CPU_Dmem_value_a5[14][2] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][30]$_SDFFE_PP0P_  (.D(net997),
    .Q(\CPU_Dmem_value_a5[14][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][31]$_SDFFE_PP0P_  (.D(net1045),
    .Q(\CPU_Dmem_value_a5[14][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][3]$_SDFFE_PP1P_  (.D(net1258),
    .Q(\CPU_Dmem_value_a5[14][3] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][4]$_SDFFE_PP0P_  (.D(net213),
    .Q(\CPU_Dmem_value_a5[14][4] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][5]$_SDFFE_PP0P_  (.D(net428),
    .Q(\CPU_Dmem_value_a5[14][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][6]$_SDFFE_PP0P_  (.D(net706),
    .Q(\CPU_Dmem_value_a5[14][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][7]$_SDFFE_PP0P_  (.D(net320),
    .Q(\CPU_Dmem_value_a5[14][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][8]$_SDFFE_PP0P_  (.D(net933),
    .Q(\CPU_Dmem_value_a5[14][8] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[14][9]$_SDFFE_PP0P_  (.D(net989),
    .Q(\CPU_Dmem_value_a5[14][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][0]$_SDFFE_PP1P_  (.D(net1205),
    .Q(\CPU_Dmem_value_a5[15][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][10]$_SDFFE_PP0P_  (.D(net732),
    .Q(\CPU_Dmem_value_a5[15][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][11]$_SDFFE_PP0P_  (.D(net306),
    .Q(\CPU_Dmem_value_a5[15][11] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][12]$_SDFFE_PP0P_  (.D(net829),
    .Q(\CPU_Dmem_value_a5[15][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][13]$_SDFFE_PP0P_  (.D(net414),
    .Q(\CPU_Dmem_value_a5[15][13] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][14]$_SDFFE_PP0P_  (.D(net312),
    .Q(\CPU_Dmem_value_a5[15][14] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][15]$_SDFFE_PP0P_  (.D(net1029),
    .Q(\CPU_Dmem_value_a5[15][15] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][16]$_SDFFE_PP0P_  (.D(net1211),
    .Q(\CPU_Dmem_value_a5[15][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][17]$_SDFFE_PP0P_  (.D(net1126),
    .Q(\CPU_Dmem_value_a5[15][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][18]$_SDFFE_PP0P_  (.D(net1100),
    .Q(\CPU_Dmem_value_a5[15][18] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][19]$_SDFFE_PP0P_  (.D(net376),
    .Q(\CPU_Dmem_value_a5[15][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][1]$_SDFFE_PP1P_  (.D(net1137),
    .Q(\CPU_Dmem_value_a5[15][1] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][20]$_SDFFE_PP0P_  (.D(net406),
    .Q(\CPU_Dmem_value_a5[15][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][21]$_SDFFE_PP0P_  (.D(net983),
    .Q(\CPU_Dmem_value_a5[15][21] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][22]$_SDFFE_PP0P_  (.D(net875),
    .Q(\CPU_Dmem_value_a5[15][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][23]$_SDFFE_PP0P_  (.D(net1025),
    .Q(\CPU_Dmem_value_a5[15][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][24]$_SDFFE_PP0P_  (.D(net294),
    .Q(\CPU_Dmem_value_a5[15][24] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][25]$_SDFFE_PP0P_  (.D(net873),
    .Q(\CPU_Dmem_value_a5[15][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][26]$_SDFFE_PP0P_  (.D(net661),
    .Q(\CPU_Dmem_value_a5[15][26] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][27]$_SDFFE_PP0P_  (.D(net426),
    .Q(\CPU_Dmem_value_a5[15][27] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][28]$_SDFFE_PP0P_  (.D(net218),
    .Q(\CPU_Dmem_value_a5[15][28] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][29]$_SDFFE_PP0P_  (.D(net971),
    .Q(\CPU_Dmem_value_a5[15][29] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][2]$_SDFFE_PP1P_  (.D(net1317),
    .Q(\CPU_Dmem_value_a5[15][2] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][30]$_SDFFE_PP0P_  (.D(net859),
    .Q(\CPU_Dmem_value_a5[15][30] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][31]$_SDFFE_PP0P_  (.D(net1133),
    .Q(\CPU_Dmem_value_a5[15][31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][3]$_SDFFE_PP1P_  (.D(net1054),
    .Q(\CPU_Dmem_value_a5[15][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][4]$_SDFFE_PP0P_  (.D(net510),
    .Q(\CPU_Dmem_value_a5[15][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][5]$_SDFFE_PP0P_  (.D(net955),
    .Q(\CPU_Dmem_value_a5[15][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][6]$_SDFFE_PP0P_  (.D(net1144),
    .Q(\CPU_Dmem_value_a5[15][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][7]$_SDFFE_PP0P_  (.D(net722),
    .Q(\CPU_Dmem_value_a5[15][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][8]$_SDFFE_PP0P_  (.D(net726),
    .Q(\CPU_Dmem_value_a5[15][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[15][9]$_SDFFE_PP0P_  (.D(net804),
    .Q(\CPU_Dmem_value_a5[15][9] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][0]$_SDFFE_PP1P_  (.D(net1115),
    .Q(\CPU_Dmem_value_a5[1][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][10]$_SDFFE_PP0P_  (.D(net613),
    .Q(\CPU_Dmem_value_a5[1][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][11]$_SDFFE_PP0P_  (.D(net927),
    .Q(\CPU_Dmem_value_a5[1][11] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][12]$_SDFFE_PP0P_  (.D(net758),
    .Q(\CPU_Dmem_value_a5[1][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][13]$_SDFFE_PP0P_  (.D(net224),
    .Q(\CPU_Dmem_value_a5[1][13] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][14]$_SDFFE_PP0P_  (.D(net262),
    .Q(\CPU_Dmem_value_a5[1][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][15]$_SDFFE_PP0P_  (.D(net734),
    .Q(\CPU_Dmem_value_a5[1][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][16]$_SDFFE_PP0P_  (.D(net392),
    .Q(\CPU_Dmem_value_a5[1][16] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][17]$_SDFFE_PP0P_  (.D(net572),
    .Q(\CPU_Dmem_value_a5[1][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][18]$_SDFFE_PP0P_  (.D(net374),
    .Q(\CPU_Dmem_value_a5[1][18] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][19]$_SDFFE_PP0P_  (.D(net1188),
    .Q(\CPU_Dmem_value_a5[1][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][1]$_SDFFE_PP0P_  (.D(net883),
    .Q(\CPU_Dmem_value_a5[1][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][20]$_SDFFE_PP0P_  (.D(net929),
    .Q(\CPU_Dmem_value_a5[1][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][21]$_SDFFE_PP0P_  (.D(net800),
    .Q(\CPU_Dmem_value_a5[1][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][22]$_SDFFE_PP0P_  (.D(net1001),
    .Q(\CPU_Dmem_value_a5[1][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][23]$_SDFFE_PP0P_  (.D(net1086),
    .Q(\CPU_Dmem_value_a5[1][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][24]$_SDFFE_PP0P_  (.D(net550),
    .Q(\CPU_Dmem_value_a5[1][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][25]$_SDFFE_PP0P_  (.D(net598),
    .Q(\CPU_Dmem_value_a5[1][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][26]$_SDFFE_PP0P_  (.D(net611),
    .Q(\CPU_Dmem_value_a5[1][26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][27]$_SDFFE_PP0P_  (.D(net390),
    .Q(\CPU_Dmem_value_a5[1][27] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][28]$_SDFFE_PP0P_  (.D(net939),
    .Q(\CPU_Dmem_value_a5[1][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][29]$_SDFFE_PP0P_  (.D(net699),
    .Q(\CPU_Dmem_value_a5[1][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][2]$_SDFFE_PP0P_  (.D(net691),
    .Q(\CPU_Dmem_value_a5[1][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][30]$_SDFFE_PP0P_  (.D(net645),
    .Q(\CPU_Dmem_value_a5[1][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][31]$_SDFFE_PP0P_  (.D(net298),
    .Q(\CPU_Dmem_value_a5[1][31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][3]$_SDFFE_PP0P_  (.D(net566),
    .Q(\CPU_Dmem_value_a5[1][3] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][4]$_SDFFE_PP0P_  (.D(net562),
    .Q(\CPU_Dmem_value_a5[1][4] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][5]$_SDFFE_PP0P_  (.D(net959),
    .Q(\CPU_Dmem_value_a5[1][5] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][6]$_SDFFE_PP0P_  (.D(net977),
    .Q(\CPU_Dmem_value_a5[1][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][7]$_SDFFE_PP0P_  (.D(net869),
    .Q(\CPU_Dmem_value_a5[1][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][8]$_SDFFE_PP0P_  (.D(net526),
    .Q(\CPU_Dmem_value_a5[1][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[1][9]$_SDFFE_PP0P_  (.D(net708),
    .Q(\CPU_Dmem_value_a5[1][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][0]$_SDFFE_PP0P_  (.D(net716),
    .Q(\CPU_Dmem_value_a5[2][0] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][10]$_SDFFE_PP0P_  (.D(net925),
    .Q(\CPU_Dmem_value_a5[2][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][11]$_SDFFE_PP0P_  (.D(net768),
    .Q(\CPU_Dmem_value_a5[2][11] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][12]$_SDFFE_PP0P_  (.D(net794),
    .Q(\CPU_Dmem_value_a5[2][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][13]$_SDFFE_PP0P_  (.D(net987),
    .Q(\CPU_Dmem_value_a5[2][13] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][14]$_SDFFE_PP0P_  (.D(net693),
    .Q(\CPU_Dmem_value_a5[2][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][15]$_SDFFE_PP0P_  (.D(net818),
    .Q(\CPU_Dmem_value_a5[2][15] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][16]$_SDFFE_PP0P_  (.D(net396),
    .Q(\CPU_Dmem_value_a5[2][16] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][17]$_SDFFE_PP0P_  (.D(net368),
    .Q(\CPU_Dmem_value_a5[2][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][18]$_SDFFE_PP0P_  (.D(net736),
    .Q(\CPU_Dmem_value_a5[2][18] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][19]$_SDFFE_PP0P_  (.D(net1011),
    .Q(\CPU_Dmem_value_a5[2][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][1]$_SDFFE_PP1P_  (.D(net1260),
    .Q(\CPU_Dmem_value_a5[2][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][20]$_SDFFE_PP0P_  (.D(net304),
    .Q(\CPU_Dmem_value_a5[2][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][21]$_SDFFE_PP0P_  (.D(net578),
    .Q(\CPU_Dmem_value_a5[2][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][22]$_SDFFE_PP0P_  (.D(net975),
    .Q(\CPU_Dmem_value_a5[2][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][23]$_SDFFE_PP0P_  (.D(net524),
    .Q(\CPU_Dmem_value_a5[2][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][24]$_SDFFE_PP0P_  (.D(net469),
    .Q(\CPU_Dmem_value_a5[2][24] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][25]$_SDFFE_PP0P_  (.D(net302),
    .Q(\CPU_Dmem_value_a5[2][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][26]$_SDFFE_PP0P_  (.D(net601),
    .Q(\CPU_Dmem_value_a5[2][26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][27]$_SDFFE_PP0P_  (.D(net398),
    .Q(\CPU_Dmem_value_a5[2][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][28]$_SDFFE_PP0P_  (.D(net704),
    .Q(\CPU_Dmem_value_a5[2][28] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][29]$_SDFFE_PP0P_  (.D(net963),
    .Q(\CPU_Dmem_value_a5[2][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][2]$_SDFFE_PP0P_  (.D(net1005),
    .Q(\CPU_Dmem_value_a5[2][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][30]$_SDFFE_PP0P_  (.D(net774),
    .Q(\CPU_Dmem_value_a5[2][30] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][31]$_SDFFE_PP0P_  (.D(net1027),
    .Q(\CPU_Dmem_value_a5[2][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][3]$_SDFFE_PP0P_  (.D(net514),
    .Q(\CPU_Dmem_value_a5[2][3] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][4]$_SDFFE_PP0P_  (.D(net485),
    .Q(\CPU_Dmem_value_a5[2][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][5]$_SDFFE_PP0P_  (.D(net1200),
    .Q(\CPU_Dmem_value_a5[2][5] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][6]$_SDFFE_PP0P_  (.D(net756),
    .Q(\CPU_Dmem_value_a5[2][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][7]$_SDFFE_PP0P_  (.D(net855),
    .Q(\CPU_Dmem_value_a5[2][7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][8]$_SDFFE_PP0P_  (.D(net280),
    .Q(\CPU_Dmem_value_a5[2][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[2][9]$_SDFFE_PP0P_  (.D(net1155),
    .Q(\CPU_Dmem_value_a5[2][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][0]$_SDFFE_PP1P_  (.D(net1414),
    .Q(\CPU_Dmem_value_a5[3][0] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][10]$_SDFFE_PP0P_  (.D(net274),
    .Q(\CPU_Dmem_value_a5[3][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][11]$_SDFFE_PP0P_  (.D(net382),
    .Q(\CPU_Dmem_value_a5[3][11] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][12]$_SDFFE_PP0P_  (.D(net326),
    .Q(\CPU_Dmem_value_a5[3][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][13]$_SDFFE_PP0P_  (.D(net677),
    .Q(\CPU_Dmem_value_a5[3][13] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][14]$_SDFFE_PP0P_  (.D(net1039),
    .Q(\CPU_Dmem_value_a5[3][14] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][15]$_SDFFE_PP0P_  (.D(net826),
    .Q(\CPU_Dmem_value_a5[3][15] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][16]$_SDFFE_PP0P_  (.D(net999),
    .Q(\CPU_Dmem_value_a5[3][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][17]$_SDFFE_PP0P_  (.D(net865),
    .Q(\CPU_Dmem_value_a5[3][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][18]$_SDFFE_PP0P_  (.D(net895),
    .Q(\CPU_Dmem_value_a5[3][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][19]$_SDFFE_PP0P_  (.D(net532),
    .Q(\CPU_Dmem_value_a5[3][19] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][1]$_SDFFE_PP1P_  (.D(net1250),
    .Q(\CPU_Dmem_value_a5[3][1] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][20]$_SDFFE_PP0P_  (.D(net238),
    .Q(\CPU_Dmem_value_a5[3][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][21]$_SDFFE_PP0P_  (.D(net278),
    .Q(\CPU_Dmem_value_a5[3][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][22]$_SDFFE_PP0P_  (.D(net1064),
    .Q(\CPU_Dmem_value_a5[3][22] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][23]$_SDFFE_PP0P_  (.D(net906),
    .Q(\CPU_Dmem_value_a5[3][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][24]$_SDFFE_PP0P_  (.D(net232),
    .Q(\CPU_Dmem_value_a5[3][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][25]$_SDFFE_PP0P_  (.D(net1021),
    .Q(\CPU_Dmem_value_a5[3][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][26]$_SDFFE_PP0P_  (.D(net290),
    .Q(\CPU_Dmem_value_a5[3][26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][27]$_SDFFE_PP0P_  (.D(net1068),
    .Q(\CPU_Dmem_value_a5[3][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][28]$_SDFFE_PP0P_  (.D(net445),
    .Q(\CPU_Dmem_value_a5[3][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][29]$_SDFFE_PP0P_  (.D(net244),
    .Q(\CPU_Dmem_value_a5[3][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][2]$_SDFFE_PP0P_  (.D(net1108),
    .Q(\CPU_Dmem_value_a5[3][2] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][30]$_SDFFE_PP0P_  (.D(net945),
    .Q(\CPU_Dmem_value_a5[3][30] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][31]$_SDFFE_PP0P_  (.D(net1117),
    .Q(\CPU_Dmem_value_a5[3][31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][3]$_SDFFE_PP0P_  (.D(net548),
    .Q(\CPU_Dmem_value_a5[3][3] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][4]$_SDFFE_PP0P_  (.D(net328),
    .Q(\CPU_Dmem_value_a5[3][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][5]$_SDFFE_PP0P_  (.D(net861),
    .Q(\CPU_Dmem_value_a5[3][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][6]$_SDFFE_PP0P_  (.D(net1165),
    .Q(\CPU_Dmem_value_a5[3][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][7]$_SDFFE_PP0P_  (.D(net1120),
    .Q(\CPU_Dmem_value_a5[3][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][8]$_SDFFE_PP0P_  (.D(net871),
    .Q(\CPU_Dmem_value_a5[3][8] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[3][9]$_SDFFE_PP0P_  (.D(net314),
    .Q(\CPU_Dmem_value_a5[3][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][0]$_SDFFE_PP0P_  (.D(net1051),
    .Q(\CPU_Dmem_value_a5[4][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][10]$_SDFFE_PP0P_  (.D(net967),
    .Q(\CPU_Dmem_value_a5[4][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][11]$_SDFFE_PP0P_  (.D(net879),
    .Q(\CPU_Dmem_value_a5[4][11] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][12]$_SDFFE_PP0P_  (.D(net1262),
    .Q(\CPU_Dmem_value_a5[4][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][13]$_SDFFE_PP0P_  (.D(net570),
    .Q(\CPU_Dmem_value_a5[4][13] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][14]$_SDFFE_PP0P_  (.D(net609),
    .Q(\CPU_Dmem_value_a5[4][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][15]$_SDFFE_PP0P_  (.D(net574),
    .Q(\CPU_Dmem_value_a5[4][15] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][16]$_SDFFE_PP0P_  (.D(net424),
    .Q(\CPU_Dmem_value_a5[4][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][17]$_SDFFE_PP0P_  (.D(net334),
    .Q(\CPU_Dmem_value_a5[4][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][18]$_SDFFE_PP0P_  (.D(net720),
    .Q(\CPU_Dmem_value_a5[4][18] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][19]$_SDFFE_PP0P_  (.D(net912),
    .Q(\CPU_Dmem_value_a5[4][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][1]$_SDFFE_PP0P_  (.D(net272),
    .Q(\CPU_Dmem_value_a5[4][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][20]$_SDFFE_PP0P_  (.D(net889),
    .Q(\CPU_Dmem_value_a5[4][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][21]$_SDFFE_PP0P_  (.D(net687),
    .Q(\CPU_Dmem_value_a5[4][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][22]$_SDFFE_PP0P_  (.D(net310),
    .Q(\CPU_Dmem_value_a5[4][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][23]$_SDFFE_PP0P_  (.D(net580),
    .Q(\CPU_Dmem_value_a5[4][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][24]$_SDFFE_PP0P_  (.D(net203),
    .Q(\CPU_Dmem_value_a5[4][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][25]$_SDFFE_PP0P_  (.D(net961),
    .Q(\CPU_Dmem_value_a5[4][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][26]$_SDFFE_PP0P_  (.D(net282),
    .Q(\CPU_Dmem_value_a5[4][26] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][27]$_SDFFE_PP0P_  (.D(net1255),
    .Q(\CPU_Dmem_value_a5[4][27] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][28]$_SDFFE_PP0P_  (.D(net808),
    .Q(\CPU_Dmem_value_a5[4][28] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][29]$_SDFFE_PP0P_  (.D(net497),
    .Q(\CPU_Dmem_value_a5[4][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][2]$_SDFFE_PP1P_  (.D(net1072),
    .Q(\CPU_Dmem_value_a5[4][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][30]$_SDFFE_PP0P_  (.D(net264),
    .Q(\CPU_Dmem_value_a5[4][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][31]$_SDFFE_PP0P_  (.D(net1070),
    .Q(\CPU_Dmem_value_a5[4][31] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][3]$_SDFFE_PP0P_  (.D(net831),
    .Q(\CPU_Dmem_value_a5[4][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][4]$_SDFFE_PP0P_  (.D(net822),
    .Q(\CPU_Dmem_value_a5[4][4] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][5]$_SDFFE_PP0P_  (.D(net1041),
    .Q(\CPU_Dmem_value_a5[4][5] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][6]$_SDFFE_PP0P_  (.D(net1159),
    .Q(\CPU_Dmem_value_a5[4][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][7]$_SDFFE_PP0P_  (.D(net760),
    .Q(\CPU_Dmem_value_a5[4][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][8]$_SDFFE_PP0P_  (.D(net487),
    .Q(\CPU_Dmem_value_a5[4][8] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[4][9]$_SDFFE_PP0P_  (.D(net1363),
    .Q(\CPU_Dmem_value_a5[4][9] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][0]$_SDFFE_PP1P_  (.D(net1314),
    .Q(\CPU_Dmem_value_a5[5][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][10]$_SDFFE_PP0P_  (.D(net1311),
    .Q(\CPU_Dmem_value_a5[5][10] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][11]$_SDFFE_PP0P_  (.D(net689),
    .Q(\CPU_Dmem_value_a5[5][11] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][12]$_SDFFE_PP0P_  (.D(net594),
    .Q(\CPU_Dmem_value_a5[5][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][13]$_SDFFE_PP0P_  (.D(net465),
    .Q(\CPU_Dmem_value_a5[5][13] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][14]$_SDFFE_PP0P_  (.D(net1181),
    .Q(\CPU_Dmem_value_a5[5][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][15]$_SDFFE_PP0P_  (.D(net354),
    .Q(\CPU_Dmem_value_a5[5][15] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][16]$_SDFFE_PP0P_  (.D(net710),
    .Q(\CPU_Dmem_value_a5[5][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][17]$_SDFFE_PP0P_  (.D(net605),
    .Q(\CPU_Dmem_value_a5[5][17] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][18]$_SDFFE_PP0P_  (.D(net495),
    .Q(\CPU_Dmem_value_a5[5][18] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][19]$_SDFFE_PP0P_  (.D(net1037),
    .Q(\CPU_Dmem_value_a5[5][19] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][1]$_SDFFE_PP0P_  (.D(net935),
    .Q(\CPU_Dmem_value_a5[5][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][20]$_SDFFE_PP0P_  (.D(net207),
    .Q(\CPU_Dmem_value_a5[5][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][21]$_SDFFE_PP0P_  (.D(net766),
    .Q(\CPU_Dmem_value_a5[5][21] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][22]$_SDFFE_PP0P_  (.D(net463),
    .Q(\CPU_Dmem_value_a5[5][22] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][23]$_SDFFE_PP0P_  (.D(net724),
    .Q(\CPU_Dmem_value_a5[5][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][24]$_SDFFE_PP0P_  (.D(net364),
    .Q(\CPU_Dmem_value_a5[5][24] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][25]$_SDFFE_PP0P_  (.D(net798),
    .Q(\CPU_Dmem_value_a5[5][25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][26]$_SDFFE_PP0P_  (.D(net916),
    .Q(\CPU_Dmem_value_a5[5][26] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][27]$_SDFFE_PP0P_  (.D(net1274),
    .Q(\CPU_Dmem_value_a5[5][27] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][28]$_SDFFE_PP0P_  (.D(net434),
    .Q(\CPU_Dmem_value_a5[5][28] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][29]$_SDFFE_PP0P_  (.D(net1003),
    .Q(\CPU_Dmem_value_a5[5][29] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][2]$_SDFFE_PP1P_  (.D(net1192),
    .Q(\CPU_Dmem_value_a5[5][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][30]$_SDFFE_PP0P_  (.D(net770),
    .Q(\CPU_Dmem_value_a5[5][30] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][31]$_SDFFE_PP0P_  (.D(net1007),
    .Q(\CPU_Dmem_value_a5[5][31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][3]$_SDFFE_PP0P_  (.D(net491),
    .Q(\CPU_Dmem_value_a5[5][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][4]$_SDFFE_PP0P_  (.D(net675),
    .Q(\CPU_Dmem_value_a5[5][4] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][5]$_SDFFE_PP0P_  (.D(net1098),
    .Q(\CPU_Dmem_value_a5[5][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][6]$_SDFFE_PP0P_  (.D(net386),
    .Q(\CPU_Dmem_value_a5[5][6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][7]$_SDFFE_PP0P_  (.D(net653),
    .Q(\CPU_Dmem_value_a5[5][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][8]$_SDFFE_PP0P_  (.D(net772),
    .Q(\CPU_Dmem_value_a5[5][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[5][9]$_SDFFE_PP0P_  (.D(net1230),
    .Q(\CPU_Dmem_value_a5[5][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][0]$_SDFFE_PP0P_  (.D(net651),
    .Q(\CPU_Dmem_value_a5[6][0] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][10]$_SDFFE_PP0P_  (.D(net340),
    .Q(\CPU_Dmem_value_a5[6][10] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][11]$_SDFFE_PP0P_  (.D(net226),
    .Q(\CPU_Dmem_value_a5[6][11] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][12]$_SDFFE_PP0P_  (.D(net270),
    .Q(\CPU_Dmem_value_a5[6][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][13]$_SDFFE_PP0P_  (.D(net1096),
    .Q(\CPU_Dmem_value_a5[6][13] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][14]$_SDFFE_PP0P_  (.D(net222),
    .Q(\CPU_Dmem_value_a5[6][14] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][15]$_SDFFE_PP0P_  (.D(net422),
    .Q(\CPU_Dmem_value_a5[6][15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][16]$_SDFFE_PP0P_  (.D(net847),
    .Q(\CPU_Dmem_value_a5[6][16] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][17]$_SDFFE_PP0P_  (.D(net346),
    .Q(\CPU_Dmem_value_a5[6][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][18]$_SDFFE_PP0P_  (.D(net332),
    .Q(\CPU_Dmem_value_a5[6][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][19]$_SDFFE_PP0P_  (.D(net619),
    .Q(\CPU_Dmem_value_a5[6][19] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][1]$_SDFFE_PP1P_  (.D(net1179),
    .Q(\CPU_Dmem_value_a5[6][1] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][20]$_SDFFE_PP0P_  (.D(net685),
    .Q(\CPU_Dmem_value_a5[6][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][21]$_SDFFE_PP0P_  (.D(net209),
    .Q(\CPU_Dmem_value_a5[6][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][22]$_SDFFE_PP0P_  (.D(net748),
    .Q(\CPU_Dmem_value_a5[6][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][23]$_SDFFE_PP0P_  (.D(net1142),
    .Q(\CPU_Dmem_value_a5[6][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][24]$_SDFFE_PP0P_  (.D(net286),
    .Q(\CPU_Dmem_value_a5[6][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][25]$_SDFFE_PP0P_  (.D(net360),
    .Q(\CPU_Dmem_value_a5[6][25] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][26]$_SDFFE_PP0P_  (.D(net669),
    .Q(\CPU_Dmem_value_a5[6][26] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][27]$_SDFFE_PP0P_  (.D(net863),
    .Q(\CPU_Dmem_value_a5[6][27] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][28]$_SDFFE_PP0P_  (.D(net416),
    .Q(\CPU_Dmem_value_a5[6][28] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][29]$_SDFFE_PP0P_  (.D(net663),
    .Q(\CPU_Dmem_value_a5[6][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][2]$_SDFFE_PP1P_  (.D(net1033),
    .Q(\CPU_Dmem_value_a5[6][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][30]$_SDFFE_PP0P_  (.D(net728),
    .Q(\CPU_Dmem_value_a5[6][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][31]$_SDFFE_PP0P_  (.D(net288),
    .Q(\CPU_Dmem_value_a5[6][31] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][3]$_SDFFE_PP0P_  (.D(net643),
    .Q(\CPU_Dmem_value_a5[6][3] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][4]$_SDFFE_PP0P_  (.D(net236),
    .Q(\CPU_Dmem_value_a5[6][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][5]$_SDFFE_PP0P_  (.D(net957),
    .Q(\CPU_Dmem_value_a5[6][5] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][6]$_SDFFE_PP0P_  (.D(net908),
    .Q(\CPU_Dmem_value_a5[6][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][7]$_SDFFE_PP0P_  (.D(net508),
    .Q(\CPU_Dmem_value_a5[6][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][8]$_SDFFE_PP0P_  (.D(net843),
    .Q(\CPU_Dmem_value_a5[6][8] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[6][9]$_SDFFE_PP0P_  (.D(net1631),
    .Q(\CPU_Dmem_value_a5[6][9] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][0]$_SDFFE_PP1P_  (.D(net1238),
    .Q(\CPU_Dmem_value_a5[7][0] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][10]$_SDFFE_PP0P_  (.D(net667),
    .Q(\CPU_Dmem_value_a5[7][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][11]$_SDFFE_PP0P_  (.D(net324),
    .Q(\CPU_Dmem_value_a5[7][11] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][12]$_SDFFE_PP0P_  (.D(net841),
    .Q(\CPU_Dmem_value_a5[7][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][13]$_SDFFE_PP0P_  (.D(net296),
    .Q(\CPU_Dmem_value_a5[7][13] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][14]$_SDFFE_PP0P_  (.D(net1066),
    .Q(\CPU_Dmem_value_a5[7][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][15]$_SDFFE_PP0P_  (.D(net584),
    .Q(\CPU_Dmem_value_a5[7][15] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][16]$_SDFFE_PP0P_  (.D(net718),
    .Q(\CPU_Dmem_value_a5[7][16] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][17]$_SDFFE_PP0P_  (.D(net623),
    .Q(\CPU_Dmem_value_a5[7][17] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][18]$_SDFFE_PP0P_  (.D(net499),
    .Q(\CPU_Dmem_value_a5[7][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][19]$_SDFFE_PP0P_  (.D(net1146),
    .Q(\CPU_Dmem_value_a5[7][19] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][1]$_SDFFE_PP1P_  (.D(net1172),
    .Q(\CPU_Dmem_value_a5[7][1] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][20]$_SDFFE_PP0P_  (.D(net308),
    .Q(\CPU_Dmem_value_a5[7][20] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][21]$_SDFFE_PP0P_  (.D(net637),
    .Q(\CPU_Dmem_value_a5[7][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][22]$_SDFFE_PP0P_  (.D(net617),
    .Q(\CPU_Dmem_value_a5[7][22] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][23]$_SDFFE_PP0P_  (.D(net1082),
    .Q(\CPU_Dmem_value_a5[7][23] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][24]$_SDFFE_PP0P_  (.D(net582),
    .Q(\CPU_Dmem_value_a5[7][24] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][25]$_SDFFE_PP0P_  (.D(net441),
    .Q(\CPU_Dmem_value_a5[7][25] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][26]$_SDFFE_PP0P_  (.D(net512),
    .Q(\CPU_Dmem_value_a5[7][26] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][27]$_SDFFE_PP0P_  (.D(net216),
    .Q(\CPU_Dmem_value_a5[7][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][28]$_SDFFE_PP0P_  (.D(net649),
    .Q(\CPU_Dmem_value_a5[7][28] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][29]$_SDFFE_PP0P_  (.D(net522),
    .Q(\CPU_Dmem_value_a5[7][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][2]$_SDFFE_PP1P_  (.D(net1080),
    .Q(\CPU_Dmem_value_a5[7][2] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][30]$_SDFFE_PP0P_  (.D(net1091),
    .Q(\CPU_Dmem_value_a5[7][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][31]$_SDFFE_PP0P_  (.D(net284),
    .Q(\CPU_Dmem_value_a5[7][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][3]$_SDFFE_PP0P_  (.D(net750),
    .Q(\CPU_Dmem_value_a5[7][3] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][4]$_SDFFE_PP0P_  (.D(net503),
    .Q(\CPU_Dmem_value_a5[7][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][5]$_SDFFE_PP0P_  (.D(net592),
    .Q(\CPU_Dmem_value_a5[7][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][6]$_SDFFE_PP0P_  (.D(net1124),
    .Q(\CPU_Dmem_value_a5[7][6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][7]$_SDFFE_PP0P_  (.D(net318),
    .Q(\CPU_Dmem_value_a5[7][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][8]$_SDFFE_PP0P_  (.D(net248),
    .Q(\CPU_Dmem_value_a5[7][8] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[7][9]$_SDFFE_PP0P_  (.D(net380),
    .Q(\CPU_Dmem_value_a5[7][9] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][0]$_SDFFE_PP0P_  (.D(net402),
    .Q(\CPU_Dmem_value_a5[8][0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][10]$_SDFFE_PP0P_  (.D(net991),
    .Q(\CPU_Dmem_value_a5[8][10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][11]$_SDFFE_PP0P_  (.D(net436),
    .Q(\CPU_Dmem_value_a5[8][11] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][12]$_SDFFE_PP0P_  (.D(net475),
    .Q(\CPU_Dmem_value_a5[8][12] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][13]$_SDFFE_PP0P_  (.D(net740),
    .Q(\CPU_Dmem_value_a5[8][13] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][14]$_SDFFE_PP0P_  (.D(net256),
    .Q(\CPU_Dmem_value_a5[8][14] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][15]$_SDFFE_PP0P_  (.D(net268),
    .Q(\CPU_Dmem_value_a5[8][15] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][16]$_SDFFE_PP0P_  (.D(net1056),
    .Q(\CPU_Dmem_value_a5[8][16] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][17]$_SDFFE_PP0P_  (.D(net322),
    .Q(\CPU_Dmem_value_a5[8][17] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][18]$_SDFFE_PP0P_  (.D(net596),
    .Q(\CPU_Dmem_value_a5[8][18] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][19]$_SDFFE_PP0P_  (.D(net449),
    .Q(\CPU_Dmem_value_a5[8][19] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][1]$_SDFFE_PP0P_  (.D(net234),
    .Q(\CPU_Dmem_value_a5[8][1] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][20]$_SDFFE_PP0P_  (.D(net639),
    .Q(\CPU_Dmem_value_a5[8][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][21]$_SDFFE_PP0P_  (.D(net404),
    .Q(\CPU_Dmem_value_a5[8][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][22]$_SDFFE_PP0P_  (.D(net744),
    .Q(\CPU_Dmem_value_a5[8][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][23]$_SDFFE_PP0P_  (.D(net919),
    .Q(\CPU_Dmem_value_a5[8][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][24]$_SDFFE_PP0P_  (.D(net937),
    .Q(\CPU_Dmem_value_a5[8][24] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][25]$_SDFFE_PP0P_  (.D(net266),
    .Q(\CPU_Dmem_value_a5[8][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][26]$_SDFFE_PP0P_  (.D(net973),
    .Q(\CPU_Dmem_value_a5[8][26] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][27]$_SDFFE_PP0P_  (.D(net853),
    .Q(\CPU_Dmem_value_a5[8][27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][28]$_SDFFE_PP0P_  (.D(net887),
    .Q(\CPU_Dmem_value_a5[8][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][29]$_SDFFE_PP0P_  (.D(net260),
    .Q(\CPU_Dmem_value_a5[8][29] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][2]$_SDFFE_PP0P_  (.D(net627),
    .Q(\CPU_Dmem_value_a5[8][2] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][30]$_SDFFE_PP0P_  (.D(net893),
    .Q(\CPU_Dmem_value_a5[8][30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][31]$_SDFFE_PP0P_  (.D(net1157),
    .Q(\CPU_Dmem_value_a5[8][31] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][3]$_SDFFE_PP1P_  (.D(net1161),
    .Q(\CPU_Dmem_value_a5[8][3] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][4]$_SDFFE_PP0P_  (.D(net338),
    .Q(\CPU_Dmem_value_a5[8][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][5]$_SDFFE_PP0P_  (.D(net1167),
    .Q(\CPU_Dmem_value_a5[8][5] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][6]$_SDFFE_PP0P_  (.D(net812),
    .Q(\CPU_Dmem_value_a5[8][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][7]$_SDFFE_PP0P_  (.D(net588),
    .Q(\CPU_Dmem_value_a5[8][7] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][8]$_SDFFE_PP0P_  (.D(net764),
    .Q(\CPU_Dmem_value_a5[8][8] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[8][9]$_SDFFE_PP0P_  (.D(net471),
    .Q(\CPU_Dmem_value_a5[8][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][0]$_SDFFE_PP1P_  (.D(net1140),
    .Q(\CPU_Dmem_value_a5[9][0] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][10]$_SDFFE_PP0P_  (.D(net1196),
    .Q(\CPU_Dmem_value_a5[9][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][11]$_SDFFE_PP0P_  (.D(net792),
    .Q(\CPU_Dmem_value_a5[9][11] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][12]$_SDFFE_PP0P_  (.D(net240),
    .Q(\CPU_Dmem_value_a5[9][12] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][13]$_SDFFE_PP0P_  (.D(net528),
    .Q(\CPU_Dmem_value_a5[9][13] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][14]$_SDFFE_PP0P_  (.D(net220),
    .Q(\CPU_Dmem_value_a5[9][14] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][15]$_SDFFE_PP0P_  (.D(net1049),
    .Q(\CPU_Dmem_value_a5[9][15] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][16]$_SDFFE_PP0P_  (.D(net246),
    .Q(\CPU_Dmem_value_a5[9][16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][17]$_SDFFE_PP0P_  (.D(net949),
    .Q(\CPU_Dmem_value_a5[9][17] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][18]$_SDFFE_PP0P_  (.D(net568),
    .Q(\CPU_Dmem_value_a5[9][18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][19]$_SDFFE_PP0P_  (.D(net564),
    .Q(\CPU_Dmem_value_a5[9][19] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][1]$_SDFFE_PP0P_  (.D(net252),
    .Q(\CPU_Dmem_value_a5[9][1] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][20]$_SDFFE_PP0P_  (.D(net205),
    .Q(\CPU_Dmem_value_a5[9][20] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][21]$_SDFFE_PP0P_  (.D(net1043),
    .Q(\CPU_Dmem_value_a5[9][21] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][22]$_SDFFE_PP0P_  (.D(net931),
    .Q(\CPU_Dmem_value_a5[9][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][23]$_SDFFE_PP0P_  (.D(net418),
    .Q(\CPU_Dmem_value_a5[9][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][24]$_SDFFE_PP0P_  (.D(net641),
    .Q(\CPU_Dmem_value_a5[9][24] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][25]$_SDFFE_PP0P_  (.D(net546),
    .Q(\CPU_Dmem_value_a5[9][25] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][26]$_SDFFE_PP0P_  (.D(net430),
    .Q(\CPU_Dmem_value_a5[9][26] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][27]$_SDFFE_PP0P_  (.D(net837),
    .Q(\CPU_Dmem_value_a5[9][27] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][28]$_SDFFE_PP0P_  (.D(net796),
    .Q(\CPU_Dmem_value_a5[9][28] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][29]$_SDFFE_PP0P_  (.D(net378),
    .Q(\CPU_Dmem_value_a5[9][29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][2]$_SDFFE_PP0P_  (.D(net1342),
    .Q(\CPU_Dmem_value_a5[9][2] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][30]$_SDFFE_PP0P_  (.D(net211),
    .Q(\CPU_Dmem_value_a5[9][30] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][31]$_SDFFE_PP0P_  (.D(net635),
    .Q(\CPU_Dmem_value_a5[9][31] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][3]$_SDFFE_PP1P_  (.D(net1322),
    .Q(\CPU_Dmem_value_a5[9][3] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][4]$_SDFFE_PP0P_  (.D(net420),
    .Q(\CPU_Dmem_value_a5[9][4] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][5]$_SDFFE_PP0P_  (.D(net833),
    .Q(\CPU_Dmem_value_a5[9][5] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][6]$_SDFFE_PP0P_  (.D(net899),
    .Q(\CPU_Dmem_value_a5[9][6] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][7]$_SDFFE_PP0P_  (.D(net536),
    .Q(\CPU_Dmem_value_a5[9][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][8]$_SDFFE_PP0P_  (.D(net659),
    .Q(\CPU_Dmem_value_a5[9][8] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Dmem_value_a5[9][9]$_SDFFE_PP0P_  (.D(net1353),
    .Q(\CPU_Dmem_value_a5[9][9] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][0]$_SDFFE_PP0P_  (.D(_00512_),
    .Q(\CPU_Xreg_value_a4[0][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][10]$_SDFFE_PP0P_  (.D(_00513_),
    .Q(\CPU_Xreg_value_a4[0][10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][11]$_SDFFE_PP0P_  (.D(_00514_),
    .Q(\CPU_Xreg_value_a4[0][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][12]$_SDFFE_PP0P_  (.D(_00515_),
    .Q(\CPU_Xreg_value_a4[0][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][13]$_SDFFE_PP0P_  (.D(_00516_),
    .Q(\CPU_Xreg_value_a4[0][13] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][14]$_SDFFE_PP0P_  (.D(_00517_),
    .Q(\CPU_Xreg_value_a4[0][14] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][15]$_SDFFE_PP0P_  (.D(_00518_),
    .Q(\CPU_Xreg_value_a4[0][15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][16]$_SDFFE_PP0P_  (.D(_00519_),
    .Q(\CPU_Xreg_value_a4[0][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][17]$_SDFFE_PP0P_  (.D(_00520_),
    .Q(\CPU_Xreg_value_a4[0][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][18]$_SDFFE_PP0P_  (.D(_00521_),
    .Q(\CPU_Xreg_value_a4[0][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][19]$_SDFFE_PP0P_  (.D(_00522_),
    .Q(\CPU_Xreg_value_a4[0][19] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][1]$_SDFFE_PP0P_  (.D(_00523_),
    .Q(\CPU_Xreg_value_a4[0][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][20]$_SDFFE_PP0P_  (.D(_00524_),
    .Q(\CPU_Xreg_value_a4[0][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][21]$_SDFFE_PP0P_  (.D(_00525_),
    .Q(\CPU_Xreg_value_a4[0][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][22]$_SDFFE_PP0P_  (.D(_00526_),
    .Q(\CPU_Xreg_value_a4[0][22] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][23]$_SDFFE_PP0P_  (.D(_00527_),
    .Q(\CPU_Xreg_value_a4[0][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][24]$_SDFFE_PP0P_  (.D(_00528_),
    .Q(\CPU_Xreg_value_a4[0][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][25]$_SDFFE_PP0P_  (.D(_00529_),
    .Q(\CPU_Xreg_value_a4[0][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][26]$_SDFFE_PP0P_  (.D(_00530_),
    .Q(\CPU_Xreg_value_a4[0][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][27]$_SDFFE_PP0P_  (.D(_00531_),
    .Q(\CPU_Xreg_value_a4[0][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][28]$_SDFFE_PP0P_  (.D(_00532_),
    .Q(\CPU_Xreg_value_a4[0][28] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][29]$_SDFFE_PP0P_  (.D(_00533_),
    .Q(\CPU_Xreg_value_a4[0][29] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][2]$_SDFFE_PP0P_  (.D(_00534_),
    .Q(\CPU_Xreg_value_a4[0][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][30]$_SDFFE_PP0P_  (.D(_00535_),
    .Q(\CPU_Xreg_value_a4[0][30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][31]$_SDFFE_PP0P_  (.D(_00536_),
    .Q(\CPU_Xreg_value_a4[0][31] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[0][3]$_SDFFE_PP0P_  (.D(_00537_),
    .Q(\CPU_Xreg_value_a4[0][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][4]$_SDFFE_PP0P_  (.D(_00538_),
    .Q(\CPU_Xreg_value_a4[0][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][5]$_SDFFE_PP0P_  (.D(_00539_),
    .Q(\CPU_Xreg_value_a4[0][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][6]$_SDFFE_PP0P_  (.D(_00540_),
    .Q(\CPU_Xreg_value_a4[0][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][7]$_SDFFE_PP0P_  (.D(_00541_),
    .Q(\CPU_Xreg_value_a4[0][7] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][8]$_SDFFE_PP0P_  (.D(_00542_),
    .Q(\CPU_Xreg_value_a4[0][8] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[0][9]$_SDFFE_PP0P_  (.D(_00543_),
    .Q(\CPU_Xreg_value_a4[0][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][0]$_SDFFE_PP0P_  (.D(_00544_),
    .Q(\CPU_Xreg_value_a4[10][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][10]$_SDFFE_PP0P_  (.D(_00545_),
    .Q(\CPU_Xreg_value_a4[10][10] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][11]$_SDFFE_PP0P_  (.D(_00546_),
    .Q(\CPU_Xreg_value_a4[10][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][12]$_SDFFE_PP0P_  (.D(_00547_),
    .Q(\CPU_Xreg_value_a4[10][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][13]$_SDFFE_PP0P_  (.D(_00548_),
    .Q(\CPU_Xreg_value_a4[10][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][14]$_SDFFE_PP0P_  (.D(_00549_),
    .Q(\CPU_Xreg_value_a4[10][14] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][15]$_SDFFE_PP0P_  (.D(_00550_),
    .Q(\CPU_Xreg_value_a4[10][15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][16]$_SDFFE_PP0P_  (.D(_00551_),
    .Q(\CPU_Xreg_value_a4[10][16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][17]$_SDFFE_PP0P_  (.D(net1574),
    .Q(\CPU_Xreg_value_a4[10][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][18]$_SDFFE_PP0P_  (.D(_00553_),
    .Q(\CPU_Xreg_value_a4[10][18] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][19]$_SDFFE_PP0P_  (.D(_00554_),
    .Q(\CPU_Xreg_value_a4[10][19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][1]$_SDFFE_PP1P_  (.D(_00555_),
    .Q(\CPU_Xreg_value_a4[10][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][20]$_SDFFE_PP0P_  (.D(net1506),
    .Q(\CPU_Xreg_value_a4[10][20] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][21]$_SDFFE_PP0P_  (.D(_00557_),
    .Q(\CPU_Xreg_value_a4[10][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][22]$_SDFFE_PP0P_  (.D(_00558_),
    .Q(\CPU_Xreg_value_a4[10][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][23]$_SDFFE_PP0P_  (.D(_00559_),
    .Q(\CPU_Xreg_value_a4[10][23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][24]$_SDFFE_PP0P_  (.D(_00560_),
    .Q(\CPU_Xreg_value_a4[10][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][25]$_SDFFE_PP0P_  (.D(_00561_),
    .Q(\CPU_Xreg_value_a4[10][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][26]$_SDFFE_PP0P_  (.D(_00562_),
    .Q(\CPU_Xreg_value_a4[10][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][27]$_SDFFE_PP0P_  (.D(_00563_),
    .Q(\CPU_Xreg_value_a4[10][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][28]$_SDFFE_PP0P_  (.D(_00564_),
    .Q(\CPU_Xreg_value_a4[10][28] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][29]$_SDFFE_PP0P_  (.D(net1563),
    .Q(\CPU_Xreg_value_a4[10][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][2]$_SDFFE_PP0P_  (.D(_00566_),
    .Q(\CPU_Xreg_value_a4[10][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][30]$_SDFFE_PP0P_  (.D(_00567_),
    .Q(\CPU_Xreg_value_a4[10][30] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][31]$_SDFFE_PP0P_  (.D(_00568_),
    .Q(\CPU_Xreg_value_a4[10][31] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][3]$_SDFFE_PP1P_  (.D(_00569_),
    .Q(\CPU_Xreg_value_a4[10][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][4]$_SDFFE_PP0P_  (.D(net1228),
    .Q(\CPU_Xreg_value_a4[10][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][5]$_SDFFE_PP0P_  (.D(_00571_),
    .Q(\CPU_Xreg_value_a4[10][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][6]$_SDFFE_PP0P_  (.D(_00572_),
    .Q(\CPU_Xreg_value_a4[10][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][7]$_SDFFE_PP0P_  (.D(_00573_),
    .Q(\CPU_Xreg_value_a4[10][7] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][8]$_SDFFE_PP0P_  (.D(_00574_),
    .Q(\CPU_Xreg_value_a4[10][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[10][9]$_SDFFE_PP0P_  (.D(_00575_),
    .Q(\CPU_Xreg_value_a4[10][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][0]$_SDFFE_PP1P_  (.D(_00576_),
    .Q(\CPU_Xreg_value_a4[11][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][10]$_SDFFE_PP0P_  (.D(_00577_),
    .Q(\CPU_Xreg_value_a4[11][10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][11]$_SDFFE_PP0P_  (.D(_00578_),
    .Q(\CPU_Xreg_value_a4[11][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][12]$_SDFFE_PP0P_  (.D(_00579_),
    .Q(\CPU_Xreg_value_a4[11][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][13]$_SDFFE_PP0P_  (.D(_00580_),
    .Q(\CPU_Xreg_value_a4[11][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][14]$_SDFFE_PP0P_  (.D(_00581_),
    .Q(\CPU_Xreg_value_a4[11][14] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][15]$_SDFFE_PP0P_  (.D(_00582_),
    .Q(\CPU_Xreg_value_a4[11][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][16]$_SDFFE_PP0P_  (.D(_00583_),
    .Q(\CPU_Xreg_value_a4[11][16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][17]$_SDFFE_PP0P_  (.D(net1532),
    .Q(\CPU_Xreg_value_a4[11][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][18]$_SDFFE_PP0P_  (.D(_00585_),
    .Q(\CPU_Xreg_value_a4[11][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][19]$_SDFFE_PP0P_  (.D(_00586_),
    .Q(\CPU_Xreg_value_a4[11][19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][1]$_SDFFE_PP1P_  (.D(_00587_),
    .Q(\CPU_Xreg_value_a4[11][1] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][20]$_SDFFE_PP0P_  (.D(_00588_),
    .Q(\CPU_Xreg_value_a4[11][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][21]$_SDFFE_PP0P_  (.D(_00589_),
    .Q(\CPU_Xreg_value_a4[11][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][22]$_SDFFE_PP0P_  (.D(_00590_),
    .Q(\CPU_Xreg_value_a4[11][22] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][23]$_SDFFE_PP0P_  (.D(_00591_),
    .Q(\CPU_Xreg_value_a4[11][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][24]$_SDFFE_PP0P_  (.D(_00592_),
    .Q(\CPU_Xreg_value_a4[11][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][25]$_SDFFE_PP0P_  (.D(_00593_),
    .Q(\CPU_Xreg_value_a4[11][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][26]$_SDFFE_PP0P_  (.D(_00594_),
    .Q(\CPU_Xreg_value_a4[11][26] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][27]$_SDFFE_PP0P_  (.D(_00595_),
    .Q(\CPU_Xreg_value_a4[11][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][28]$_SDFFE_PP0P_  (.D(_00596_),
    .Q(\CPU_Xreg_value_a4[11][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][29]$_SDFFE_PP0P_  (.D(_00597_),
    .Q(\CPU_Xreg_value_a4[11][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][2]$_SDFFE_PP0P_  (.D(_00598_),
    .Q(\CPU_Xreg_value_a4[11][2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][30]$_SDFFE_PP0P_  (.D(_00599_),
    .Q(\CPU_Xreg_value_a4[11][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][31]$_SDFFE_PP0P_  (.D(_00600_),
    .Q(\CPU_Xreg_value_a4[11][31] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][3]$_SDFFE_PP1P_  (.D(_00601_),
    .Q(\CPU_Xreg_value_a4[11][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][4]$_SDFFE_PP0P_  (.D(net1218),
    .Q(\CPU_Xreg_value_a4[11][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][5]$_SDFFE_PP0P_  (.D(_00603_),
    .Q(\CPU_Xreg_value_a4[11][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][6]$_SDFFE_PP0P_  (.D(_00604_),
    .Q(\CPU_Xreg_value_a4[11][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][7]$_SDFFE_PP0P_  (.D(_00605_),
    .Q(\CPU_Xreg_value_a4[11][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][8]$_SDFFE_PP0P_  (.D(_00606_),
    .Q(\CPU_Xreg_value_a4[11][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[11][9]$_SDFFE_PP0P_  (.D(_00607_),
    .Q(\CPU_Xreg_value_a4[11][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][0]$_SDFFE_PP0P_  (.D(_00608_),
    .Q(\CPU_Xreg_value_a4[12][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][10]$_SDFFE_PP0P_  (.D(_00609_),
    .Q(\CPU_Xreg_value_a4[12][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][11]$_SDFFE_PP0P_  (.D(_00610_),
    .Q(\CPU_Xreg_value_a4[12][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][12]$_SDFFE_PP0P_  (.D(_00611_),
    .Q(\CPU_Xreg_value_a4[12][12] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][13]$_SDFFE_PP0P_  (.D(_00612_),
    .Q(\CPU_Xreg_value_a4[12][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][14]$_SDFFE_PP0P_  (.D(_00613_),
    .Q(\CPU_Xreg_value_a4[12][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][15]$_SDFFE_PP0P_  (.D(_00614_),
    .Q(\CPU_Xreg_value_a4[12][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][16]$_SDFFE_PP0P_  (.D(_00615_),
    .Q(\CPU_Xreg_value_a4[12][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][17]$_SDFFE_PP0P_  (.D(net1567),
    .Q(\CPU_Xreg_value_a4[12][17] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][18]$_SDFFE_PP0P_  (.D(_00617_),
    .Q(\CPU_Xreg_value_a4[12][18] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][19]$_SDFFE_PP0P_  (.D(_00618_),
    .Q(\CPU_Xreg_value_a4[12][19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][1]$_SDFFE_PP0P_  (.D(_00619_),
    .Q(\CPU_Xreg_value_a4[12][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][20]$_SDFFE_PP0P_  (.D(_00620_),
    .Q(\CPU_Xreg_value_a4[12][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][21]$_SDFFE_PP0P_  (.D(_00621_),
    .Q(\CPU_Xreg_value_a4[12][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][22]$_SDFFE_PP0P_  (.D(_00622_),
    .Q(\CPU_Xreg_value_a4[12][22] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][23]$_SDFFE_PP0P_  (.D(_00623_),
    .Q(\CPU_Xreg_value_a4[12][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][24]$_SDFFE_PP0P_  (.D(_00624_),
    .Q(\CPU_Xreg_value_a4[12][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][25]$_SDFFE_PP0P_  (.D(_00625_),
    .Q(\CPU_Xreg_value_a4[12][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][26]$_SDFFE_PP0P_  (.D(_00626_),
    .Q(\CPU_Xreg_value_a4[12][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][27]$_SDFFE_PP0P_  (.D(_00627_),
    .Q(\CPU_Xreg_value_a4[12][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][28]$_SDFFE_PP0P_  (.D(_00628_),
    .Q(\CPU_Xreg_value_a4[12][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][29]$_SDFFE_PP0P_  (.D(_00629_),
    .Q(\CPU_Xreg_value_a4[12][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][2]$_SDFFE_PP1P_  (.D(_00630_),
    .Q(\CPU_Xreg_value_a4[12][2] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][30]$_SDFFE_PP0P_  (.D(_00631_),
    .Q(\CPU_Xreg_value_a4[12][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][31]$_SDFFE_PP0P_  (.D(_00632_),
    .Q(\CPU_Xreg_value_a4[12][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][3]$_SDFFE_PP1P_  (.D(_00633_),
    .Q(\CPU_Xreg_value_a4[12][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][4]$_SDFFE_PP0P_  (.D(net1286),
    .Q(\CPU_Xreg_value_a4[12][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][5]$_SDFFE_PP0P_  (.D(_00635_),
    .Q(\CPU_Xreg_value_a4[12][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][6]$_SDFFE_PP0P_  (.D(_00636_),
    .Q(\CPU_Xreg_value_a4[12][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][7]$_SDFFE_PP0P_  (.D(_00637_),
    .Q(\CPU_Xreg_value_a4[12][7] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][8]$_SDFFE_PP0P_  (.D(_00638_),
    .Q(\CPU_Xreg_value_a4[12][8] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[12][9]$_SDFFE_PP0P_  (.D(_00639_),
    .Q(\CPU_Xreg_value_a4[12][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][0]$_SDFFE_PP1P_  (.D(_00640_),
    .Q(\CPU_Xreg_value_a4[13][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][10]$_SDFFE_PP0P_  (.D(_00641_),
    .Q(\CPU_Xreg_value_a4[13][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][11]$_SDFFE_PP0P_  (.D(_00642_),
    .Q(\CPU_Xreg_value_a4[13][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][12]$_SDFFE_PP0P_  (.D(_00643_),
    .Q(\CPU_Xreg_value_a4[13][12] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][13]$_SDFFE_PP0P_  (.D(_00644_),
    .Q(\CPU_Xreg_value_a4[13][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][14]$_SDFFE_PP0P_  (.D(_00645_),
    .Q(\CPU_Xreg_value_a4[13][14] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][15]$_SDFFE_PP0P_  (.D(_00646_),
    .Q(\CPU_Xreg_value_a4[13][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][16]$_SDFFE_PP0P_  (.D(_00647_),
    .Q(\CPU_Xreg_value_a4[13][16] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][17]$_SDFFE_PP0P_  (.D(net1603),
    .Q(\CPU_Xreg_value_a4[13][17] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][18]$_SDFFE_PP0P_  (.D(_00649_),
    .Q(\CPU_Xreg_value_a4[13][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][19]$_SDFFE_PP0P_  (.D(_00650_),
    .Q(\CPU_Xreg_value_a4[13][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][1]$_SDFFE_PP0P_  (.D(_00651_),
    .Q(\CPU_Xreg_value_a4[13][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][20]$_SDFFE_PP0P_  (.D(net1648),
    .Q(\CPU_Xreg_value_a4[13][20] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][21]$_SDFFE_PP0P_  (.D(_00653_),
    .Q(\CPU_Xreg_value_a4[13][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][22]$_SDFFE_PP0P_  (.D(_00654_),
    .Q(\CPU_Xreg_value_a4[13][22] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][23]$_SDFFE_PP0P_  (.D(_00655_),
    .Q(\CPU_Xreg_value_a4[13][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][24]$_SDFFE_PP0P_  (.D(_00656_),
    .Q(\CPU_Xreg_value_a4[13][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][25]$_SDFFE_PP0P_  (.D(_00657_),
    .Q(\CPU_Xreg_value_a4[13][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][26]$_SDFFE_PP0P_  (.D(_00658_),
    .Q(\CPU_Xreg_value_a4[13][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][27]$_SDFFE_PP0P_  (.D(_00659_),
    .Q(\CPU_Xreg_value_a4[13][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][28]$_SDFFE_PP0P_  (.D(_00660_),
    .Q(\CPU_Xreg_value_a4[13][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][29]$_SDFFE_PP0P_  (.D(net1536),
    .Q(\CPU_Xreg_value_a4[13][29] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][2]$_SDFFE_PP1P_  (.D(_00662_),
    .Q(\CPU_Xreg_value_a4[13][2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][30]$_SDFFE_PP0P_  (.D(_00663_),
    .Q(\CPU_Xreg_value_a4[13][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][31]$_SDFFE_PP0P_  (.D(_00664_),
    .Q(\CPU_Xreg_value_a4[13][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][3]$_SDFFE_PP1P_  (.D(_00665_),
    .Q(\CPU_Xreg_value_a4[13][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][4]$_SDFFE_PP0P_  (.D(net1198),
    .Q(\CPU_Xreg_value_a4[13][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][5]$_SDFFE_PP0P_  (.D(_00667_),
    .Q(\CPU_Xreg_value_a4[13][5] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][6]$_SDFFE_PP0P_  (.D(_00668_),
    .Q(\CPU_Xreg_value_a4[13][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][7]$_SDFFE_PP0P_  (.D(_00669_),
    .Q(\CPU_Xreg_value_a4[13][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][8]$_SDFFE_PP0P_  (.D(_00670_),
    .Q(\CPU_Xreg_value_a4[13][8] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[13][9]$_SDFFE_PP0P_  (.D(_00671_),
    .Q(\CPU_Xreg_value_a4[13][9] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[14][0]$_SDFFE_PP0P_  (.D(_00672_),
    .Q(\CPU_Xreg_value_a4[14][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][10]$_SDFFE_PP0P_  (.D(_00673_),
    .Q(\CPU_Xreg_value_a4[14][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][11]$_SDFFE_PP0P_  (.D(_00674_),
    .Q(\CPU_Xreg_value_a4[14][11] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][12]$_SDFFE_PP0P_  (.D(_00675_),
    .Q(\CPU_Xreg_value_a4[14][12] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][13]$_SDFFE_PP0P_  (.D(_00676_),
    .Q(\CPU_Xreg_value_a4[14][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][14]$_SDFFE_PP0P_  (.D(_00677_),
    .Q(\CPU_Xreg_value_a4[14][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][15]$_SDFFE_PP0P_  (.D(_00678_),
    .Q(\CPU_Xreg_value_a4[14][15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][16]$_SDFFE_PP0P_  (.D(_00679_),
    .Q(\CPU_Xreg_value_a4[14][16] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][17]$_SDFFE_PP0P_  (.D(net1513),
    .Q(\CPU_Xreg_value_a4[14][17] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][18]$_SDFFE_PP0P_  (.D(_00681_),
    .Q(\CPU_Xreg_value_a4[14][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][19]$_SDFFE_PP0P_  (.D(_00682_),
    .Q(\CPU_Xreg_value_a4[14][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][1]$_SDFFE_PP1P_  (.D(_00683_),
    .Q(\CPU_Xreg_value_a4[14][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][20]$_SDFFE_PP0P_  (.D(net1592),
    .Q(\CPU_Xreg_value_a4[14][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][21]$_SDFFE_PP0P_  (.D(_00685_),
    .Q(\CPU_Xreg_value_a4[14][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][22]$_SDFFE_PP0P_  (.D(_00686_),
    .Q(\CPU_Xreg_value_a4[14][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][23]$_SDFFE_PP0P_  (.D(_00687_),
    .Q(\CPU_Xreg_value_a4[14][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][24]$_SDFFE_PP0P_  (.D(_00688_),
    .Q(\CPU_Xreg_value_a4[14][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][25]$_SDFFE_PP0P_  (.D(_00689_),
    .Q(\CPU_Xreg_value_a4[14][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][26]$_SDFFE_PP0P_  (.D(_00690_),
    .Q(\CPU_Xreg_value_a4[14][26] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][27]$_SDFFE_PP0P_  (.D(_00691_),
    .Q(\CPU_Xreg_value_a4[14][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][28]$_SDFFE_PP0P_  (.D(_00692_),
    .Q(\CPU_Xreg_value_a4[14][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][29]$_SDFFE_PP0P_  (.D(net1560),
    .Q(\CPU_Xreg_value_a4[14][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][2]$_SDFFE_PP1P_  (.D(_00694_),
    .Q(\CPU_Xreg_value_a4[14][2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][30]$_SDFFE_PP0P_  (.D(_00695_),
    .Q(\CPU_Xreg_value_a4[14][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][31]$_SDFFE_PP0P_  (.D(_00696_),
    .Q(\CPU_Xreg_value_a4[14][31] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][3]$_SDFFE_PP1P_  (.D(_00697_),
    .Q(\CPU_Xreg_value_a4[14][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][4]$_SDFFE_PP0P_  (.D(_00698_),
    .Q(\CPU_Xreg_value_a4[14][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[14][5]$_SDFFE_PP0P_  (.D(_00699_),
    .Q(\CPU_Xreg_value_a4[14][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][6]$_SDFFE_PP0P_  (.D(_00700_),
    .Q(\CPU_Xreg_value_a4[14][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[14][7]$_SDFFE_PP0P_  (.D(_00701_),
    .Q(\CPU_Xreg_value_a4[14][7] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[14][8]$_SDFFE_PP0P_  (.D(_00702_),
    .Q(\CPU_Xreg_value_a4[14][8] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_Xreg_value_a4[14][9]$_SDFFE_PP0P_  (.D(_00703_),
    .Q(\CPU_Xreg_value_a4[14][9] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][0]$_SDFFE_PP1P_  (.D(_00704_),
    .Q(\CPU_Xreg_value_a4[15][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][10]$_SDFFE_PP0P_  (.D(_00705_),
    .Q(\CPU_Xreg_value_a4[15][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][11]$_SDFFE_PP0P_  (.D(_00706_),
    .Q(\CPU_Xreg_value_a4[15][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][12]$_SDFFE_PP0P_  (.D(_00707_),
    .Q(\CPU_Xreg_value_a4[15][12] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][13]$_SDFFE_PP0P_  (.D(_00708_),
    .Q(\CPU_Xreg_value_a4[15][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][14]$_SDFFE_PP0P_  (.D(_00709_),
    .Q(\CPU_Xreg_value_a4[15][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][15]$_SDFFE_PP0P_  (.D(_00710_),
    .Q(\CPU_Xreg_value_a4[15][15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][16]$_SDFFE_PP0P_  (.D(_00711_),
    .Q(\CPU_Xreg_value_a4[15][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][17]$_SDFFE_PP0P_  (.D(net1499),
    .Q(\CPU_Xreg_value_a4[15][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][18]$_SDFFE_PP0P_  (.D(_00713_),
    .Q(\CPU_Xreg_value_a4[15][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][19]$_SDFFE_PP0P_  (.D(_00714_),
    .Q(\CPU_Xreg_value_a4[15][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][1]$_SDFFE_PP1P_  (.D(_00715_),
    .Q(\CPU_Xreg_value_a4[15][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][20]$_SDFFE_PP0P_  (.D(net1654),
    .Q(\CPU_Xreg_value_a4[15][20] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][21]$_SDFFE_PP0P_  (.D(_00717_),
    .Q(\CPU_Xreg_value_a4[15][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][22]$_SDFFE_PP0P_  (.D(_00718_),
    .Q(\CPU_Xreg_value_a4[15][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][23]$_SDFFE_PP0P_  (.D(_00719_),
    .Q(\CPU_Xreg_value_a4[15][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][24]$_SDFFE_PP0P_  (.D(_00720_),
    .Q(\CPU_Xreg_value_a4[15][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][25]$_SDFFE_PP0P_  (.D(_00721_),
    .Q(\CPU_Xreg_value_a4[15][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][26]$_SDFFE_PP0P_  (.D(_00722_),
    .Q(\CPU_Xreg_value_a4[15][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][27]$_SDFFE_PP0P_  (.D(_00723_),
    .Q(\CPU_Xreg_value_a4[15][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][28]$_SDFFE_PP0P_  (.D(_00724_),
    .Q(\CPU_Xreg_value_a4[15][28] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][29]$_SDFFE_PP0P_  (.D(net1594),
    .Q(\CPU_Xreg_value_a4[15][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][2]$_SDFFE_PP1P_  (.D(_00726_),
    .Q(\CPU_Xreg_value_a4[15][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][30]$_SDFFE_PP0P_  (.D(_00727_),
    .Q(\CPU_Xreg_value_a4[15][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][31]$_SDFFE_PP0P_  (.D(_00728_),
    .Q(\CPU_Xreg_value_a4[15][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][3]$_SDFFE_PP1P_  (.D(_00729_),
    .Q(\CPU_Xreg_value_a4[15][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][4]$_SDFFE_PP0P_  (.D(net1272),
    .Q(\CPU_Xreg_value_a4[15][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][5]$_SDFFE_PP0P_  (.D(_00731_),
    .Q(\CPU_Xreg_value_a4[15][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][6]$_SDFFE_PP0P_  (.D(_00732_),
    .Q(\CPU_Xreg_value_a4[15][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][7]$_SDFFE_PP0P_  (.D(_00733_),
    .Q(\CPU_Xreg_value_a4[15][7] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][8]$_SDFFE_PP0P_  (.D(_00734_),
    .Q(\CPU_Xreg_value_a4[15][8] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[15][9]$_SDFFE_PP0P_  (.D(_00735_),
    .Q(\CPU_Xreg_value_a4[15][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][0]$_SDFFE_PP1P_  (.D(_00736_),
    .Q(\CPU_Xreg_value_a4[1][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][10]$_SDFFE_PP0P_  (.D(_00737_),
    .Q(\CPU_Xreg_value_a4[1][10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][11]$_SDFFE_PP0P_  (.D(_00738_),
    .Q(\CPU_Xreg_value_a4[1][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][12]$_SDFFE_PP0P_  (.D(_00739_),
    .Q(\CPU_Xreg_value_a4[1][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][13]$_SDFFE_PP0P_  (.D(_00740_),
    .Q(\CPU_Xreg_value_a4[1][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][14]$_SDFFE_PP0P_  (.D(_00741_),
    .Q(\CPU_Xreg_value_a4[1][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][15]$_SDFFE_PP0P_  (.D(_00742_),
    .Q(\CPU_Xreg_value_a4[1][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][16]$_SDFFE_PP0P_  (.D(_00743_),
    .Q(\CPU_Xreg_value_a4[1][16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][17]$_SDFFE_PP0P_  (.D(net1645),
    .Q(\CPU_Xreg_value_a4[1][17] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][18]$_SDFFE_PP0P_  (.D(_00745_),
    .Q(\CPU_Xreg_value_a4[1][18] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][19]$_SDFFE_PP0P_  (.D(_00746_),
    .Q(\CPU_Xreg_value_a4[1][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][1]$_SDFFE_PP0P_  (.D(_00747_),
    .Q(\CPU_Xreg_value_a4[1][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][20]$_SDFFE_PP0P_  (.D(net1587),
    .Q(\CPU_Xreg_value_a4[1][20] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][21]$_SDFFE_PP0P_  (.D(_00749_),
    .Q(\CPU_Xreg_value_a4[1][21] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][22]$_SDFFE_PP0P_  (.D(_00750_),
    .Q(\CPU_Xreg_value_a4[1][22] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][23]$_SDFFE_PP0P_  (.D(_00751_),
    .Q(\CPU_Xreg_value_a4[1][23] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][24]$_SDFFE_PP0P_  (.D(_00752_),
    .Q(\CPU_Xreg_value_a4[1][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][25]$_SDFFE_PP0P_  (.D(_00753_),
    .Q(\CPU_Xreg_value_a4[1][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][26]$_SDFFE_PP0P_  (.D(_00754_),
    .Q(\CPU_Xreg_value_a4[1][26] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][27]$_SDFFE_PP0P_  (.D(_00755_),
    .Q(\CPU_Xreg_value_a4[1][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][28]$_SDFFE_PP0P_  (.D(_00756_),
    .Q(\CPU_Xreg_value_a4[1][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][29]$_SDFFE_PP0P_  (.D(net1634),
    .Q(\CPU_Xreg_value_a4[1][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][2]$_SDFFE_PP0P_  (.D(_00758_),
    .Q(\CPU_Xreg_value_a4[1][2] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][30]$_SDFFE_PP0P_  (.D(_00759_),
    .Q(\CPU_Xreg_value_a4[1][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][31]$_SDFFE_PP0P_  (.D(_00760_),
    .Q(\CPU_Xreg_value_a4[1][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][3]$_SDFFE_PP0P_  (.D(_00761_),
    .Q(\CPU_Xreg_value_a4[1][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][4]$_SDFFE_PP0P_  (.D(net1281),
    .Q(\CPU_Xreg_value_a4[1][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][5]$_SDFFE_PP0P_  (.D(_00763_),
    .Q(\CPU_Xreg_value_a4[1][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][6]$_SDFFE_PP0P_  (.D(_00764_),
    .Q(\CPU_Xreg_value_a4[1][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][7]$_SDFFE_PP0P_  (.D(_00765_),
    .Q(\CPU_Xreg_value_a4[1][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][8]$_SDFFE_PP0P_  (.D(_00766_),
    .Q(\CPU_Xreg_value_a4[1][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[1][9]$_SDFFE_PP0P_  (.D(_00767_),
    .Q(\CPU_Xreg_value_a4[1][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][0]$_SDFFE_PP0P_  (.D(_00768_),
    .Q(\CPU_Xreg_value_a4[2][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][10]$_SDFFE_PP0P_  (.D(_00769_),
    .Q(\CPU_Xreg_value_a4[2][10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][11]$_SDFFE_PP0P_  (.D(_00770_),
    .Q(\CPU_Xreg_value_a4[2][11] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][12]$_SDFFE_PP0P_  (.D(_00771_),
    .Q(\CPU_Xreg_value_a4[2][12] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][13]$_SDFFE_PP0P_  (.D(_00772_),
    .Q(\CPU_Xreg_value_a4[2][13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][14]$_SDFFE_PP0P_  (.D(_00773_),
    .Q(\CPU_Xreg_value_a4[2][14] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][15]$_SDFFE_PP0P_  (.D(_00774_),
    .Q(\CPU_Xreg_value_a4[2][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][16]$_SDFFE_PP0P_  (.D(_00775_),
    .Q(\CPU_Xreg_value_a4[2][16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][17]$_SDFFE_PP0P_  (.D(net1642),
    .Q(\CPU_Xreg_value_a4[2][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][18]$_SDFFE_PP0P_  (.D(_00777_),
    .Q(\CPU_Xreg_value_a4[2][18] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][19]$_SDFFE_PP0P_  (.D(_00778_),
    .Q(\CPU_Xreg_value_a4[2][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][1]$_SDFFE_PP1P_  (.D(_00779_),
    .Q(\CPU_Xreg_value_a4[2][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][20]$_SDFFE_PP0P_  (.D(_00780_),
    .Q(\CPU_Xreg_value_a4[2][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][21]$_SDFFE_PP0P_  (.D(_00781_),
    .Q(\CPU_Xreg_value_a4[2][21] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][22]$_SDFFE_PP0P_  (.D(_00782_),
    .Q(\CPU_Xreg_value_a4[2][22] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][23]$_SDFFE_PP0P_  (.D(_00783_),
    .Q(\CPU_Xreg_value_a4[2][23] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][24]$_SDFFE_PP0P_  (.D(_00784_),
    .Q(\CPU_Xreg_value_a4[2][24] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][25]$_SDFFE_PP0P_  (.D(_00785_),
    .Q(\CPU_Xreg_value_a4[2][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][26]$_SDFFE_PP0P_  (.D(_00786_),
    .Q(\CPU_Xreg_value_a4[2][26] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][27]$_SDFFE_PP0P_  (.D(_00787_),
    .Q(\CPU_Xreg_value_a4[2][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][28]$_SDFFE_PP0P_  (.D(_00788_),
    .Q(\CPU_Xreg_value_a4[2][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][29]$_SDFFE_PP0P_  (.D(_00789_),
    .Q(\CPU_Xreg_value_a4[2][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][2]$_SDFFE_PP0P_  (.D(_00790_),
    .Q(\CPU_Xreg_value_a4[2][2] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][30]$_SDFFE_PP0P_  (.D(_00791_),
    .Q(\CPU_Xreg_value_a4[2][30] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][31]$_SDFFE_PP0P_  (.D(_00792_),
    .Q(\CPU_Xreg_value_a4[2][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][3]$_SDFFE_PP0P_  (.D(_00793_),
    .Q(\CPU_Xreg_value_a4[2][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][4]$_SDFFE_PP0P_  (.D(net1277),
    .Q(\CPU_Xreg_value_a4[2][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][5]$_SDFFE_PP0P_  (.D(_00795_),
    .Q(\CPU_Xreg_value_a4[2][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][6]$_SDFFE_PP0P_  (.D(_00796_),
    .Q(\CPU_Xreg_value_a4[2][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][7]$_SDFFE_PP0P_  (.D(_00797_),
    .Q(\CPU_Xreg_value_a4[2][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][8]$_SDFFE_PP0P_  (.D(_00798_),
    .Q(\CPU_Xreg_value_a4[2][8] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[2][9]$_SDFFE_PP0P_  (.D(_00799_),
    .Q(\CPU_Xreg_value_a4[2][9] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][0]$_SDFFE_PP1P_  (.D(_00800_),
    .Q(\CPU_Xreg_value_a4[3][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][10]$_SDFFE_PP0P_  (.D(_00801_),
    .Q(\CPU_Xreg_value_a4[3][10] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][11]$_SDFFE_PP0P_  (.D(_00802_),
    .Q(\CPU_Xreg_value_a4[3][11] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][12]$_SDFFE_PP0P_  (.D(_00803_),
    .Q(\CPU_Xreg_value_a4[3][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][13]$_SDFFE_PP0P_  (.D(_00804_),
    .Q(\CPU_Xreg_value_a4[3][13] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][14]$_SDFFE_PP0P_  (.D(_00805_),
    .Q(\CPU_Xreg_value_a4[3][14] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][15]$_SDFFE_PP0P_  (.D(_00806_),
    .Q(\CPU_Xreg_value_a4[3][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][16]$_SDFFE_PP0P_  (.D(_00807_),
    .Q(\CPU_Xreg_value_a4[3][16] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][17]$_SDFFE_PP0P_  (.D(net1550),
    .Q(\CPU_Xreg_value_a4[3][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][18]$_SDFFE_PP0P_  (.D(_00809_),
    .Q(\CPU_Xreg_value_a4[3][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][19]$_SDFFE_PP0P_  (.D(_00810_),
    .Q(\CPU_Xreg_value_a4[3][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][1]$_SDFFE_PP1P_  (.D(_00811_),
    .Q(\CPU_Xreg_value_a4[3][1] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][20]$_SDFFE_PP0P_  (.D(_00812_),
    .Q(\CPU_Xreg_value_a4[3][20] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][21]$_SDFFE_PP0P_  (.D(_00813_),
    .Q(\CPU_Xreg_value_a4[3][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][22]$_SDFFE_PP0P_  (.D(_00814_),
    .Q(\CPU_Xreg_value_a4[3][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][23]$_SDFFE_PP0P_  (.D(_00815_),
    .Q(\CPU_Xreg_value_a4[3][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][24]$_SDFFE_PP0P_  (.D(_00816_),
    .Q(\CPU_Xreg_value_a4[3][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][25]$_SDFFE_PP0P_  (.D(_00817_),
    .Q(\CPU_Xreg_value_a4[3][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][26]$_SDFFE_PP0P_  (.D(_00818_),
    .Q(\CPU_Xreg_value_a4[3][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][27]$_SDFFE_PP0P_  (.D(_00819_),
    .Q(\CPU_Xreg_value_a4[3][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][28]$_SDFFE_PP0P_  (.D(_00820_),
    .Q(\CPU_Xreg_value_a4[3][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][29]$_SDFFE_PP0P_  (.D(net1638),
    .Q(\CPU_Xreg_value_a4[3][29] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][2]$_SDFFE_PP0P_  (.D(_00822_),
    .Q(\CPU_Xreg_value_a4[3][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][30]$_SDFFE_PP0P_  (.D(_00823_),
    .Q(\CPU_Xreg_value_a4[3][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][31]$_SDFFE_PP0P_  (.D(_00824_),
    .Q(\CPU_Xreg_value_a4[3][31] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][3]$_SDFFE_PP0P_  (.D(_00825_),
    .Q(\CPU_Xreg_value_a4[3][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][4]$_SDFFE_PP0P_  (.D(net1183),
    .Q(\CPU_Xreg_value_a4[3][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][5]$_SDFFE_PP0P_  (.D(_00827_),
    .Q(\CPU_Xreg_value_a4[3][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][6]$_SDFFE_PP0P_  (.D(_00828_),
    .Q(\CPU_Xreg_value_a4[3][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][7]$_SDFFE_PP0P_  (.D(_00829_),
    .Q(\CPU_Xreg_value_a4[3][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][8]$_SDFFE_PP0P_  (.D(_00830_),
    .Q(\CPU_Xreg_value_a4[3][8] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[3][9]$_SDFFE_PP0P_  (.D(_00831_),
    .Q(\CPU_Xreg_value_a4[3][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][0]$_SDFFE_PP0P_  (.D(_00832_),
    .Q(\CPU_Xreg_value_a4[4][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][10]$_SDFFE_PP0P_  (.D(_00833_),
    .Q(\CPU_Xreg_value_a4[4][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][11]$_SDFFE_PP0P_  (.D(_00834_),
    .Q(\CPU_Xreg_value_a4[4][11] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][12]$_SDFFE_PP0P_  (.D(_00835_),
    .Q(\CPU_Xreg_value_a4[4][12] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][13]$_SDFFE_PP0P_  (.D(_00836_),
    .Q(\CPU_Xreg_value_a4[4][13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][14]$_SDFFE_PP0P_  (.D(_00837_),
    .Q(\CPU_Xreg_value_a4[4][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][15]$_SDFFE_PP0P_  (.D(_00838_),
    .Q(\CPU_Xreg_value_a4[4][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][16]$_SDFFE_PP0P_  (.D(_00839_),
    .Q(\CPU_Xreg_value_a4[4][16] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][17]$_SDFFE_PP0P_  (.D(net1527),
    .Q(\CPU_Xreg_value_a4[4][17] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][18]$_SDFFE_PP0P_  (.D(_00841_),
    .Q(\CPU_Xreg_value_a4[4][18] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][19]$_SDFFE_PP0P_  (.D(_00842_),
    .Q(\CPU_Xreg_value_a4[4][19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][1]$_SDFFE_PP0P_  (.D(_00843_),
    .Q(\CPU_Xreg_value_a4[4][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][20]$_SDFFE_PP0P_  (.D(_00844_),
    .Q(\CPU_Xreg_value_a4[4][20] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][21]$_SDFFE_PP0P_  (.D(_00845_),
    .Q(\CPU_Xreg_value_a4[4][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][22]$_SDFFE_PP0P_  (.D(_00846_),
    .Q(\CPU_Xreg_value_a4[4][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][23]$_SDFFE_PP0P_  (.D(_00847_),
    .Q(\CPU_Xreg_value_a4[4][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][24]$_SDFFE_PP0P_  (.D(_00848_),
    .Q(\CPU_Xreg_value_a4[4][24] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][25]$_SDFFE_PP0P_  (.D(_00849_),
    .Q(\CPU_Xreg_value_a4[4][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][26]$_SDFFE_PP0P_  (.D(_00850_),
    .Q(\CPU_Xreg_value_a4[4][26] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][27]$_SDFFE_PP0P_  (.D(_00851_),
    .Q(\CPU_Xreg_value_a4[4][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][28]$_SDFFE_PP0P_  (.D(_00852_),
    .Q(\CPU_Xreg_value_a4[4][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][29]$_SDFFE_PP0P_  (.D(_00853_),
    .Q(\CPU_Xreg_value_a4[4][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][2]$_SDFFE_PP1P_  (.D(_00854_),
    .Q(\CPU_Xreg_value_a4[4][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][30]$_SDFFE_PP0P_  (.D(_00855_),
    .Q(\CPU_Xreg_value_a4[4][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][31]$_SDFFE_PP0P_  (.D(_00856_),
    .Q(\CPU_Xreg_value_a4[4][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][3]$_SDFFE_PP0P_  (.D(_00857_),
    .Q(\CPU_Xreg_value_a4[4][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][4]$_SDFFE_PP0P_  (.D(net1169),
    .Q(\CPU_Xreg_value_a4[4][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][5]$_SDFFE_PP0P_  (.D(_00859_),
    .Q(\CPU_Xreg_value_a4[4][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][6]$_SDFFE_PP0P_  (.D(_00860_),
    .Q(\CPU_Xreg_value_a4[4][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][7]$_SDFFE_PP0P_  (.D(_00861_),
    .Q(\CPU_Xreg_value_a4[4][7] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][8]$_SDFFE_PP0P_  (.D(_00862_),
    .Q(\CPU_Xreg_value_a4[4][8] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[4][9]$_SDFFE_PP0P_  (.D(_00863_),
    .Q(\CPU_Xreg_value_a4[4][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][0]$_SDFFE_PP1P_  (.D(_00864_),
    .Q(\CPU_Xreg_value_a4[5][0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][10]$_SDFFE_PP0P_  (.D(_00865_),
    .Q(\CPU_Xreg_value_a4[5][10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][11]$_SDFFE_PP0P_  (.D(_00866_),
    .Q(\CPU_Xreg_value_a4[5][11] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][12]$_SDFFE_PP0P_  (.D(_00867_),
    .Q(\CPU_Xreg_value_a4[5][12] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][13]$_SDFFE_PP0P_  (.D(_00868_),
    .Q(\CPU_Xreg_value_a4[5][13] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][14]$_SDFFE_PP0P_  (.D(_00869_),
    .Q(\CPU_Xreg_value_a4[5][14] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][15]$_SDFFE_PP0P_  (.D(_00870_),
    .Q(\CPU_Xreg_value_a4[5][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][16]$_SDFFE_PP0P_  (.D(_00871_),
    .Q(\CPU_Xreg_value_a4[5][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][17]$_SDFFE_PP0P_  (.D(net1606),
    .Q(\CPU_Xreg_value_a4[5][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][18]$_SDFFE_PP0P_  (.D(_00873_),
    .Q(\CPU_Xreg_value_a4[5][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][19]$_SDFFE_PP0P_  (.D(_00874_),
    .Q(\CPU_Xreg_value_a4[5][19] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][1]$_SDFFE_PP0P_  (.D(_00875_),
    .Q(\CPU_Xreg_value_a4[5][1] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][20]$_SDFFE_PP0P_  (.D(net1525),
    .Q(\CPU_Xreg_value_a4[5][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][21]$_SDFFE_PP0P_  (.D(_00877_),
    .Q(\CPU_Xreg_value_a4[5][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][22]$_SDFFE_PP0P_  (.D(_00878_),
    .Q(\CPU_Xreg_value_a4[5][22] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][23]$_SDFFE_PP0P_  (.D(_00879_),
    .Q(\CPU_Xreg_value_a4[5][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][24]$_SDFFE_PP0P_  (.D(_00880_),
    .Q(\CPU_Xreg_value_a4[5][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][25]$_SDFFE_PP0P_  (.D(_00881_),
    .Q(\CPU_Xreg_value_a4[5][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][26]$_SDFFE_PP0P_  (.D(_00882_),
    .Q(\CPU_Xreg_value_a4[5][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][27]$_SDFFE_PP0P_  (.D(_00883_),
    .Q(\CPU_Xreg_value_a4[5][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][28]$_SDFFE_PP0P_  (.D(_00884_),
    .Q(\CPU_Xreg_value_a4[5][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][29]$_SDFFE_PP0P_  (.D(net1620),
    .Q(\CPU_Xreg_value_a4[5][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][2]$_SDFFE_PP1P_  (.D(_00886_),
    .Q(\CPU_Xreg_value_a4[5][2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][30]$_SDFFE_PP0P_  (.D(_00887_),
    .Q(\CPU_Xreg_value_a4[5][30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][31]$_SDFFE_PP0P_  (.D(_00888_),
    .Q(\CPU_Xreg_value_a4[5][31] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][3]$_SDFFE_PP0P_  (.D(_00889_),
    .Q(\CPU_Xreg_value_a4[5][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][4]$_SDFFE_PP0P_  (.D(net1240),
    .Q(\CPU_Xreg_value_a4[5][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][5]$_SDFFE_PP0P_  (.D(_00891_),
    .Q(\CPU_Xreg_value_a4[5][5] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][6]$_SDFFE_PP0P_  (.D(_00892_),
    .Q(\CPU_Xreg_value_a4[5][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][7]$_SDFFE_PP0P_  (.D(_00893_),
    .Q(\CPU_Xreg_value_a4[5][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][8]$_SDFFE_PP0P_  (.D(_00894_),
    .Q(\CPU_Xreg_value_a4[5][8] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[5][9]$_SDFFE_PP0P_  (.D(_00895_),
    .Q(\CPU_Xreg_value_a4[5][9] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][0]$_SDFFE_PP0P_  (.D(_00896_),
    .Q(\CPU_Xreg_value_a4[6][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][10]$_SDFFE_PP0P_  (.D(_00897_),
    .Q(\CPU_Xreg_value_a4[6][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][11]$_SDFFE_PP0P_  (.D(_00898_),
    .Q(\CPU_Xreg_value_a4[6][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][12]$_SDFFE_PP0P_  (.D(_00899_),
    .Q(\CPU_Xreg_value_a4[6][12] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][13]$_SDFFE_PP0P_  (.D(_00900_),
    .Q(\CPU_Xreg_value_a4[6][13] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][14]$_SDFFE_PP0P_  (.D(_00901_),
    .Q(\CPU_Xreg_value_a4[6][14] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][15]$_SDFFE_PP0P_  (.D(_00902_),
    .Q(\CPU_Xreg_value_a4[6][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][16]$_SDFFE_PP0P_  (.D(_00903_),
    .Q(\CPU_Xreg_value_a4[6][16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][17]$_SDFFE_PP0P_  (.D(net1661),
    .Q(\CPU_Xreg_value_a4[6][17] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][18]$_SDFFE_PP0P_  (.D(_00905_),
    .Q(\CPU_Xreg_value_a4[6][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][19]$_SDFFE_PP0P_  (.D(_00906_),
    .Q(\CPU_Xreg_value_a4[6][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][1]$_SDFFE_PP1P_  (.D(_00907_),
    .Q(\CPU_Xreg_value_a4[6][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][20]$_SDFFE_PP0P_  (.D(_00908_),
    .Q(\CPU_Xreg_value_a4[6][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][21]$_SDFFE_PP0P_  (.D(_00909_),
    .Q(\CPU_Xreg_value_a4[6][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][22]$_SDFFE_PP0P_  (.D(_00910_),
    .Q(\CPU_Xreg_value_a4[6][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][23]$_SDFFE_PP0P_  (.D(_00911_),
    .Q(\CPU_Xreg_value_a4[6][23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][24]$_SDFFE_PP0P_  (.D(_00912_),
    .Q(\CPU_Xreg_value_a4[6][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][25]$_SDFFE_PP0P_  (.D(_00913_),
    .Q(\CPU_Xreg_value_a4[6][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][26]$_SDFFE_PP0P_  (.D(_00914_),
    .Q(\CPU_Xreg_value_a4[6][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][27]$_SDFFE_PP0P_  (.D(_00915_),
    .Q(\CPU_Xreg_value_a4[6][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][28]$_SDFFE_PP0P_  (.D(_00916_),
    .Q(\CPU_Xreg_value_a4[6][28] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][29]$_SDFFE_PP0P_  (.D(_00917_),
    .Q(\CPU_Xreg_value_a4[6][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][2]$_SDFFE_PP1P_  (.D(_00918_),
    .Q(\CPU_Xreg_value_a4[6][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][30]$_SDFFE_PP0P_  (.D(_00919_),
    .Q(\CPU_Xreg_value_a4[6][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][31]$_SDFFE_PP0P_  (.D(_00920_),
    .Q(\CPU_Xreg_value_a4[6][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][3]$_SDFFE_PP0P_  (.D(_00921_),
    .Q(\CPU_Xreg_value_a4[6][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][4]$_SDFFE_PP0P_  (.D(net1244),
    .Q(\CPU_Xreg_value_a4[6][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][5]$_SDFFE_PP0P_  (.D(_00923_),
    .Q(\CPU_Xreg_value_a4[6][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][6]$_SDFFE_PP0P_  (.D(_00924_),
    .Q(\CPU_Xreg_value_a4[6][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][7]$_SDFFE_PP0P_  (.D(_00925_),
    .Q(\CPU_Xreg_value_a4[6][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][8]$_SDFFE_PP0P_  (.D(_00926_),
    .Q(\CPU_Xreg_value_a4[6][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[6][9]$_SDFFE_PP0P_  (.D(_00927_),
    .Q(\CPU_Xreg_value_a4[6][9] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][0]$_SDFFE_PP1P_  (.D(_00928_),
    .Q(\CPU_Xreg_value_a4[7][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][10]$_SDFFE_PP0P_  (.D(_00929_),
    .Q(\CPU_Xreg_value_a4[7][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][11]$_SDFFE_PP0P_  (.D(_00930_),
    .Q(\CPU_Xreg_value_a4[7][11] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][12]$_SDFFE_PP0P_  (.D(_00931_),
    .Q(\CPU_Xreg_value_a4[7][12] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][13]$_SDFFE_PP0P_  (.D(_00932_),
    .Q(\CPU_Xreg_value_a4[7][13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][14]$_SDFFE_PP0P_  (.D(_00933_),
    .Q(\CPU_Xreg_value_a4[7][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][15]$_SDFFE_PP0P_  (.D(_00934_),
    .Q(\CPU_Xreg_value_a4[7][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][16]$_SDFFE_PP0P_  (.D(_00935_),
    .Q(\CPU_Xreg_value_a4[7][16] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][17]$_SDFFE_PP0P_  (.D(net1578),
    .Q(\CPU_Xreg_value_a4[7][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][18]$_SDFFE_PP0P_  (.D(_00937_),
    .Q(\CPU_Xreg_value_a4[7][18] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][19]$_SDFFE_PP0P_  (.D(_00938_),
    .Q(\CPU_Xreg_value_a4[7][19] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][1]$_SDFFE_PP1P_  (.D(_00939_),
    .Q(\CPU_Xreg_value_a4[7][1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][20]$_SDFFE_PP0P_  (.D(_00940_),
    .Q(\CPU_Xreg_value_a4[7][20] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][21]$_SDFFE_PP0P_  (.D(_00941_),
    .Q(\CPU_Xreg_value_a4[7][21] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][22]$_SDFFE_PP0P_  (.D(_00942_),
    .Q(\CPU_Xreg_value_a4[7][22] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][23]$_SDFFE_PP0P_  (.D(_00943_),
    .Q(\CPU_Xreg_value_a4[7][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][24]$_SDFFE_PP0P_  (.D(_00944_),
    .Q(\CPU_Xreg_value_a4[7][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][25]$_SDFFE_PP0P_  (.D(_00945_),
    .Q(\CPU_Xreg_value_a4[7][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][26]$_SDFFE_PP0P_  (.D(_00946_),
    .Q(\CPU_Xreg_value_a4[7][26] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][27]$_SDFFE_PP0P_  (.D(_00947_),
    .Q(\CPU_Xreg_value_a4[7][27] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][28]$_SDFFE_PP0P_  (.D(_00948_),
    .Q(\CPU_Xreg_value_a4[7][28] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][29]$_SDFFE_PP0P_  (.D(net1509),
    .Q(\CPU_Xreg_value_a4[7][29] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][2]$_SDFFE_PP1P_  (.D(_00950_),
    .Q(\CPU_Xreg_value_a4[7][2] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][30]$_SDFFE_PP0P_  (.D(_00951_),
    .Q(\CPU_Xreg_value_a4[7][30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][31]$_SDFFE_PP0P_  (.D(_00952_),
    .Q(\CPU_Xreg_value_a4[7][31] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][3]$_SDFFE_PP0P_  (.D(_00953_),
    .Q(\CPU_Xreg_value_a4[7][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][4]$_SDFFE_PP0P_  (.D(net1339),
    .Q(\CPU_Xreg_value_a4[7][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][5]$_SDFFE_PP0P_  (.D(_00955_),
    .Q(\CPU_Xreg_value_a4[7][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][6]$_SDFFE_PP0P_  (.D(_00956_),
    .Q(\CPU_Xreg_value_a4[7][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][7]$_SDFFE_PP0P_  (.D(_00957_),
    .Q(\CPU_Xreg_value_a4[7][7] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][8]$_SDFFE_PP0P_  (.D(_00958_),
    .Q(\CPU_Xreg_value_a4[7][8] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[7][9]$_SDFFE_PP0P_  (.D(_00959_),
    .Q(\CPU_Xreg_value_a4[7][9] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][0]$_SDFFE_PP0P_  (.D(_00960_),
    .Q(\CPU_Xreg_value_a4[8][0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][10]$_SDFFE_PP0P_  (.D(_00961_),
    .Q(\CPU_Xreg_value_a4[8][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][11]$_SDFFE_PP0P_  (.D(_00962_),
    .Q(\CPU_Xreg_value_a4[8][11] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][12]$_SDFFE_PP0P_  (.D(_00963_),
    .Q(\CPU_Xreg_value_a4[8][12] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][13]$_SDFFE_PP0P_  (.D(_00964_),
    .Q(\CPU_Xreg_value_a4[8][13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][14]$_SDFFE_PP0P_  (.D(_00965_),
    .Q(\CPU_Xreg_value_a4[8][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][15]$_SDFFE_PP0P_  (.D(_00966_),
    .Q(\CPU_Xreg_value_a4[8][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][16]$_SDFFE_PP0P_  (.D(_00967_),
    .Q(\CPU_Xreg_value_a4[8][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][17]$_SDFFE_PP0P_  (.D(net1596),
    .Q(\CPU_Xreg_value_a4[8][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][18]$_SDFFE_PP0P_  (.D(_00969_),
    .Q(\CPU_Xreg_value_a4[8][18] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][19]$_SDFFE_PP0P_  (.D(_00970_),
    .Q(\CPU_Xreg_value_a4[8][19] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][1]$_SDFFE_PP0P_  (.D(_00971_),
    .Q(\CPU_Xreg_value_a4[8][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][20]$_SDFFE_PP0P_  (.D(_00972_),
    .Q(\CPU_Xreg_value_a4[8][20] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][21]$_SDFFE_PP0P_  (.D(_00973_),
    .Q(\CPU_Xreg_value_a4[8][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][22]$_SDFFE_PP0P_  (.D(_00974_),
    .Q(\CPU_Xreg_value_a4[8][22] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][23]$_SDFFE_PP0P_  (.D(_00975_),
    .Q(\CPU_Xreg_value_a4[8][23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][24]$_SDFFE_PP0P_  (.D(_00976_),
    .Q(\CPU_Xreg_value_a4[8][24] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][25]$_SDFFE_PP0P_  (.D(_00977_),
    .Q(\CPU_Xreg_value_a4[8][25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][26]$_SDFFE_PP0P_  (.D(_00978_),
    .Q(\CPU_Xreg_value_a4[8][26] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][27]$_SDFFE_PP0P_  (.D(_00979_),
    .Q(\CPU_Xreg_value_a4[8][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][28]$_SDFFE_PP0P_  (.D(_00980_),
    .Q(\CPU_Xreg_value_a4[8][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][29]$_SDFFE_PP0P_  (.D(net1548),
    .Q(\CPU_Xreg_value_a4[8][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][2]$_SDFFE_PP0P_  (.D(_00982_),
    .Q(\CPU_Xreg_value_a4[8][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][30]$_SDFFE_PP0P_  (.D(_00983_),
    .Q(\CPU_Xreg_value_a4[8][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][31]$_SDFFE_PP0P_  (.D(_00984_),
    .Q(\CPU_Xreg_value_a4[8][31] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][3]$_SDFFE_PP1P_  (.D(_00985_),
    .Q(\CPU_Xreg_value_a4[8][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][4]$_SDFFE_PP0P_  (.D(net1150),
    .Q(\CPU_Xreg_value_a4[8][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][5]$_SDFFE_PP0P_  (.D(_00987_),
    .Q(\CPU_Xreg_value_a4[8][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][6]$_SDFFE_PP0P_  (.D(_00988_),
    .Q(\CPU_Xreg_value_a4[8][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][7]$_SDFFE_PP0P_  (.D(_00989_),
    .Q(\CPU_Xreg_value_a4[8][7] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][8]$_SDFFE_PP0P_  (.D(_00990_),
    .Q(\CPU_Xreg_value_a4[8][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[8][9]$_SDFFE_PP0P_  (.D(_00991_),
    .Q(\CPU_Xreg_value_a4[8][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][0]$_SDFFE_PP1P_  (.D(_00992_),
    .Q(\CPU_Xreg_value_a4[9][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][10]$_SDFFE_PP0P_  (.D(_00993_),
    .Q(\CPU_Xreg_value_a4[9][10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][11]$_SDFFE_PP0P_  (.D(_00994_),
    .Q(\CPU_Xreg_value_a4[9][11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][12]$_SDFFE_PP0P_  (.D(_00995_),
    .Q(\CPU_Xreg_value_a4[9][12] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][13]$_SDFFE_PP0P_  (.D(_00996_),
    .Q(\CPU_Xreg_value_a4[9][13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][14]$_SDFFE_PP0P_  (.D(_00997_),
    .Q(\CPU_Xreg_value_a4[9][14] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][15]$_SDFFE_PP0P_  (.D(_00998_),
    .Q(\CPU_Xreg_value_a4[9][15] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][16]$_SDFFE_PP0P_  (.D(_00999_),
    .Q(\CPU_Xreg_value_a4[9][16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][17]$_SDFFE_PP0P_  (.D(net1544),
    .Q(\CPU_Xreg_value_a4[9][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][18]$_SDFFE_PP0P_  (.D(_01001_),
    .Q(\CPU_Xreg_value_a4[9][18] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][19]$_SDFFE_PP0P_  (.D(_01002_),
    .Q(\CPU_Xreg_value_a4[9][19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][1]$_SDFFE_PP0P_  (.D(_01003_),
    .Q(\CPU_Xreg_value_a4[9][1] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][20]$_SDFFE_PP0P_  (.D(net1657),
    .Q(\CPU_Xreg_value_a4[9][20] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][21]$_SDFFE_PP0P_  (.D(_01005_),
    .Q(\CPU_Xreg_value_a4[9][21] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][22]$_SDFFE_PP0P_  (.D(_01006_),
    .Q(\CPU_Xreg_value_a4[9][22] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][23]$_SDFFE_PP0P_  (.D(_01007_),
    .Q(\CPU_Xreg_value_a4[9][23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][24]$_SDFFE_PP0P_  (.D(_01008_),
    .Q(\CPU_Xreg_value_a4[9][24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][25]$_SDFFE_PP0P_  (.D(_01009_),
    .Q(\CPU_Xreg_value_a4[9][25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][26]$_SDFFE_PP0P_  (.D(_01010_),
    .Q(\CPU_Xreg_value_a4[9][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][27]$_SDFFE_PP0P_  (.D(_01011_),
    .Q(\CPU_Xreg_value_a4[9][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][28]$_SDFFE_PP0P_  (.D(_01012_),
    .Q(\CPU_Xreg_value_a4[9][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][29]$_SDFFE_PP0P_  (.D(net1529),
    .Q(\CPU_Xreg_value_a4[9][29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][2]$_SDFFE_PP0P_  (.D(_01014_),
    .Q(\CPU_Xreg_value_a4[9][2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][30]$_SDFFE_PP0P_  (.D(_01015_),
    .Q(\CPU_Xreg_value_a4[9][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][31]$_SDFFE_PP0P_  (.D(_01016_),
    .Q(\CPU_Xreg_value_a4[9][31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][3]$_SDFFE_PP1P_  (.D(_01017_),
    .Q(\CPU_Xreg_value_a4[9][3] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][4]$_SDFFE_PP0P_  (.D(net1328),
    .Q(\CPU_Xreg_value_a4[9][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][5]$_SDFFE_PP0P_  (.D(_01019_),
    .Q(\CPU_Xreg_value_a4[9][5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][6]$_SDFFE_PP0P_  (.D(_01020_),
    .Q(\CPU_Xreg_value_a4[9][6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][7]$_SDFFE_PP0P_  (.D(_01021_),
    .Q(\CPU_Xreg_value_a4[9][7] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][8]$_SDFFE_PP0P_  (.D(_01022_),
    .Q(\CPU_Xreg_value_a4[9][8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a4[9][9]$_SDFFE_PP0P_  (.D(_01023_),
    .Q(\CPU_Xreg_value_a4[9][9] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][0]$_DFF_P_  (.D(net191),
    .Q(\CPU_Xreg_value_a5[14][0] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][1]$_DFF_P_  (.D(net171),
    .Q(\CPU_Xreg_value_a5[14][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][2]$_DFF_P_  (.D(net168),
    .Q(\CPU_Xreg_value_a5[14][2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][3]$_DFF_P_  (.D(net186),
    .Q(\CPU_Xreg_value_a5[14][3] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][4]$_DFF_P_  (.D(net166),
    .Q(\CPU_Xreg_value_a5[14][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][5]$_DFF_P_  (.D(net180),
    .Q(\CPU_Xreg_value_a5[14][5] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][6]$_DFF_P_  (.D(net165),
    .Q(\CPU_Xreg_value_a5[14][6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][7]$_DFF_P_  (.D(net504),
    .Q(\CPU_Xreg_value_a5[14][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][8]$_DFF_P_  (.D(net195),
    .Q(\CPU_Xreg_value_a5[14][8] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_Xreg_value_a5[14][9]$_DFF_P_  (.D(net172),
    .Q(\CPU_Xreg_value_a5[14][9] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[0]$_DFF_P_  (.D(\CPU_br_tgt_pc_a2[0] ),
    .Q(\CPU_br_tgt_pc_a3[0] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[1]$_DFF_P_  (.D(\CPU_br_tgt_pc_a2[1] ),
    .Q(\CPU_br_tgt_pc_a3[1] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[2]$_DFF_P_  (.D(\CPU_br_tgt_pc_a2[2] ),
    .Q(\CPU_br_tgt_pc_a3[2] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[3]$_DFF_P_  (.D(\CPU_br_tgt_pc_a2[3] ),
    .Q(\CPU_br_tgt_pc_a3[3] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[4]$_DFF_P_  (.D(net1716),
    .Q(\CPU_br_tgt_pc_a3[4] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_br_tgt_pc_a3[5]$_DFF_P_  (.D(net1694),
    .Q(\CPU_br_tgt_pc_a3[5] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[0]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[0] ),
    .Q(\CPU_dmem_rd_data_a5[0] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[10]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[10] ),
    .Q(\CPU_dmem_rd_data_a5[10] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[11]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[11] ),
    .Q(\CPU_dmem_rd_data_a5[11] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[12]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[12] ),
    .Q(\CPU_dmem_rd_data_a5[12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[13]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[13] ),
    .Q(\CPU_dmem_rd_data_a5[13] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[14]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[14] ),
    .Q(\CPU_dmem_rd_data_a5[14] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[15]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[15] ),
    .Q(\CPU_dmem_rd_data_a5[15] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[16]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[16] ),
    .Q(\CPU_dmem_rd_data_a5[16] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[17]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[17] ),
    .Q(\CPU_dmem_rd_data_a5[17] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[18]$_DFF_P_  (.D(net1789),
    .Q(\CPU_dmem_rd_data_a5[18] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[19]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[19] ),
    .Q(\CPU_dmem_rd_data_a5[19] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[1]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[1] ),
    .Q(\CPU_dmem_rd_data_a5[1] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[20]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[20] ),
    .Q(\CPU_dmem_rd_data_a5[20] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[21]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[21] ),
    .Q(\CPU_dmem_rd_data_a5[21] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[22]$_DFF_P_  (.D(net1755),
    .Q(\CPU_dmem_rd_data_a5[22] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_dmem_rd_data_a5[23]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[23] ),
    .Q(\CPU_dmem_rd_data_a5[23] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[24]$_DFF_P_  (.D(net1709),
    .Q(\CPU_dmem_rd_data_a5[24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[25]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[25] ),
    .Q(\CPU_dmem_rd_data_a5[25] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[26]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[26] ),
    .Q(\CPU_dmem_rd_data_a5[26] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[27]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[27] ),
    .Q(\CPU_dmem_rd_data_a5[27] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[28]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[28] ),
    .Q(\CPU_dmem_rd_data_a5[28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[29]$_DFF_P_  (.D(net1822),
    .Q(\CPU_dmem_rd_data_a5[29] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[2]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[2] ),
    .Q(\CPU_dmem_rd_data_a5[2] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[30]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[30] ),
    .Q(\CPU_dmem_rd_data_a5[30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[31]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[31] ),
    .Q(\CPU_dmem_rd_data_a5[31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[3]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[3] ),
    .Q(\CPU_dmem_rd_data_a5[3] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[4]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[4] ),
    .Q(\CPU_dmem_rd_data_a5[4] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[5]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[5] ),
    .Q(\CPU_dmem_rd_data_a5[5] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[6]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[6] ),
    .Q(\CPU_dmem_rd_data_a5[6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[7]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[7] ),
    .Q(\CPU_dmem_rd_data_a5[7] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_dmem_rd_data_a5[8]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[8] ),
    .Q(\CPU_dmem_rd_data_a5[8] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_dmem_rd_data_a5[9]$_DFF_P_  (.D(\w_CPU_dmem_rd_data_a4[9] ),
    .Q(\CPU_dmem_rd_data_a5[9] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_imem_rd_addr_a1[0]$_SDFF_PP0_  (.D(_01024_),
    .Q(\CPU_imem_rd_addr_a1[0] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_imem_rd_addr_a1[1]$_SDFF_PP0_  (.D(net1017),
    .Q(\CPU_imem_rd_addr_a1[1] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_imem_rd_addr_a1[2]$_SDFF_PP0_  (.D(net1558),
    .Q(\CPU_imem_rd_addr_a1[2] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_imem_rd_addr_a1[3]$_SDFF_PP0_  (.D(net1583),
    .Q(\CPU_imem_rd_addr_a1[3] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[0]$_DFF_P_  (.D(\CPU_imm_a1[0] ),
    .Q(\CPU_imm_a2[0] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[11]$_DFF_P_  (.D(\CPU_imm_a1[11] ),
    .Q(\CPU_imm_a2[11] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[1]$_DFF_P_  (.D(\CPU_imm_a1[1] ),
    .Q(\CPU_imm_a2[1] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[2]$_DFF_P_  (.D(\CPU_imm_a1[2] ),
    .Q(\CPU_imm_a2[2] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[30]$_DFF_P_  (.D(\CPU_imm_a1[10] ),
    .Q(\CPU_imm_a2[10] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[3]$_DFF_P_  (.D(\CPU_imm_a1[3] ),
    .Q(\CPU_imm_a2[3] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a2[4]$_SDFF_PP0_  (.D(_01028_),
    .Q(\CPU_imm_a2[4] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a3[0]$_DFF_P_  (.D(net150),
    .Q(\CPU_imm_a3[0] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_imm_a3[11]$_DFF_P_  (.D(net145),
    .Q(\CPU_imm_a3[11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a3[1]$_DFF_P_  (.D(net159),
    .Q(\CPU_imm_a3[1] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a3[2]$_DFF_P_  (.D(net161),
    .Q(\CPU_imm_a3[2] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_imm_a3[30]$_DFF_P_  (.D(net179),
    .Q(\CPU_imm_a3[10] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a3[3]$_DFF_P_  (.D(net155),
    .Q(\CPU_imm_a3[3] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_imm_a3[4]$_DFF_P_  (.D(net152),
    .Q(\CPU_imm_a3[4] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[0]$_DFF_P_  (.D(net138),
    .Q(\CPU_inc_pc_a2[0] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[1]$_DFF_P_  (.D(net148),
    .Q(\CPU_inc_pc_a2[1] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[2]$_DFF_P_  (.D(\CPU_inc_pc_a1[2] ),
    .Q(\CPU_inc_pc_a2[2] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[3]$_DFF_P_  (.D(\CPU_inc_pc_a1[3] ),
    .Q(\CPU_inc_pc_a2[3] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[4]$_DFF_P_  (.D(\CPU_inc_pc_a1[4] ),
    .Q(\CPU_inc_pc_a2[4] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a2[5]$_DFF_P_  (.D(\CPU_inc_pc_a1[5] ),
    .Q(\CPU_inc_pc_a2[5] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[0]$_DFF_P_  (.D(net154),
    .Q(\CPU_inc_pc_a3[0] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[1]$_DFF_P_  (.D(net156),
    .Q(\CPU_inc_pc_a3[1] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[2]$_DFF_P_  (.D(net129),
    .Q(\CPU_inc_pc_a3[2] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[3]$_DFF_P_  (.D(net128),
    .Q(\CPU_inc_pc_a3[3] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[4]$_DFF_P_  (.D(net123),
    .Q(\CPU_inc_pc_a3[4] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_inc_pc_a3[5]$_DFF_P_  (.D(net124),
    .Q(\CPU_inc_pc_a3[5] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_add_a2$_DFF_P_  (.D(CPU_is_add_a1),
    .Q(CPU_is_add_a2),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_is_add_a3$_DFF_P_  (.D(net139),
    .Q(CPU_is_add_a3),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_addi_a2$_DFF_P_  (.D(CPU_is_addi_a1),
    .Q(CPU_is_addi_a2),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_is_addi_a3$_DFF_P_  (.D(net118),
    .Q(CPU_is_addi_a3),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_blt_a2$_DFF_P_  (.D(CPU_is_blt_a1),
    .Q(CPU_is_blt_a2),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_blt_a3$_DFF_P_  (.D(net133),
    .Q(CPU_is_blt_a3),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_bltu_a2$_DFF_P_  (.D(net111),
    .Q(CPU_is_bltu_a2),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_bltu_a3$_DFF_P_  (.D(net146),
    .Q(CPU_is_bltu_a3),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_load_a2$_DFF_P_  (.D(CPU_is_load_a1),
    .Q(CPU_is_load_a2),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_load_a3$_DFF_P_  (.D(net116),
    .Q(CPU_is_load_a3),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_s_instr_a2$_DFF_P_  (.D(CPU_is_s_instr_a1),
    .Q(CPU_is_s_instr_a2),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_s_instr_a3$_DFF_P_  (.D(net131),
    .Q(CPU_is_s_instr_a3),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_is_s_instr_a4$_DFF_P_  (.D(net115),
    .Q(CPU_is_s_instr_a4),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_slt_a2$_DFF_P_  (.D(net112),
    .Q(CPU_is_slt_a2),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_slt_a3$_DFF_P_  (.D(net141),
    .Q(CPU_is_slt_a3),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_slti_a2$_DFF_P_  (.D(net113),
    .Q(CPU_is_slti_a2),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_is_slti_a3$_DFF_P_  (.D(net149),
    .Q(CPU_is_slti_a3),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a1[0]$_SDFFE_PP0P_  (.D(net752),
    .Q(\CPU_inc_pc_a1[0] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a1[1]$_SDFFE_PP0P_  (.D(net1031),
    .Q(\CPU_inc_pc_a1[1] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a2[2]$_DFF_P_  (.D(net192),
    .Q(\CPU_pc_a2[2] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a2[3]$_DFF_P_  (.D(net182),
    .Q(\CPU_pc_a2[3] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a2[4]$_DFF_P_  (.D(net827),
    .Q(\CPU_pc_a2[4] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_pc_a2[5]$_DFF_P_  (.D(net1291),
    .Q(\CPU_pc_a2[5] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a2[0]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[7] ),
    .Q(\CPU_rd_a2[0] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a2[1]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[8] ),
    .Q(\CPU_rd_a2[1] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a2[2]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[9] ),
    .Q(\CPU_rd_a2[2] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a2[3]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[10] ),
    .Q(\CPU_rd_a2[3] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a2[4]$_DFF_P_  (.D(\CPU_dec_bits_a1[10] ),
    .Q(\CPU_rd_a2[4] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_rd_a3[0]$_DFF_P_  (.D(net121),
    .Q(\CPU_rd_a3[0] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_rd_a3[1]$_DFF_P_  (.D(net117),
    .Q(\CPU_rd_a3[1] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rd_a3[2]$_DFF_P_  (.D(net130),
    .Q(\CPU_rd_a3[2] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rd_a3[3]$_DFF_P_  (.D(net119),
    .Q(\CPU_rd_a3[3] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_rd_a3[4]$_DFF_P_  (.D(net136),
    .Q(\CPU_rd_a3[4] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a4[0]$_DFF_P_  (.D(net177),
    .Q(\CPU_rd_a4[0] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a4[1]$_DFF_P_  (.D(net900),
    .Q(\CPU_rd_a4[1] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a4[2]$_DFF_P_  (.D(net1104),
    .Q(\CPU_rd_a4[2] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a4[3]$_DFF_P_  (.D(net1263),
    .Q(\CPU_rd_a4[3] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a4[4]$_DFF_P_  (.D(net174),
    .Q(\CPU_rd_a4[4] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a5[0]$_DFF_P_  (.D(net127),
    .Q(\CPU_rd_a5[0] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a5[1]$_DFF_P_  (.D(net114),
    .Q(\CPU_rd_a5[1] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a5[2]$_DFF_P_  (.D(net125),
    .Q(\CPU_rd_a5[2] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a5[3]$_DFF_P_  (.D(net122),
    .Q(\CPU_rd_a5[3] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_a5[4]$_DFF_P_  (.D(net126),
    .Q(\CPU_rd_a5[4] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_valid_a2$_DFF_P_  (.D(CPU_rd_valid_a1),
    .Q(CPU_rd_valid_a2),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_rd_valid_a3$_DFF_P_  (.D(net132),
    .Q(CPU_rd_valid_a3),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_reset_a1$_DFF_P_  (.D(net1),
    .Q(CPU_reset_a1),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_reset_a2$_DFF_P_  (.D(net1214),
    .Q(CPU_reset_a2),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_reset_a3$_DFF_P_  (.D(net120),
    .Q(CPU_reset_a3),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_reset_a4$_DFF_P_  (.D(net108),
    .Q(CPU_reset_a4),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_result_a4[0]$_DFF_P_  (.D(\CPU_result_a3[2] ),
    .Q(\CPU_dmem_addr_a4[0] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_result_a4[1]$_DFF_P_  (.D(\CPU_result_a3[3] ),
    .Q(\CPU_dmem_addr_a4[1] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_result_a4[2]$_DFF_P_  (.D(\CPU_result_a3[4] ),
    .Q(\CPU_dmem_addr_a4[2] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_result_a4[3]$_DFF_P_  (.D(\CPU_result_a3[5] ),
    .Q(\CPU_dmem_addr_a4[3] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs1_a2[0]$_SDFF_PN0_  (.D(_01031_),
    .Q(\CPU_rf_rd_index1_a2[0] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs1_a2[1]$_SDFF_PN0_  (.D(_01032_),
    .Q(\CPU_rf_rd_index1_a2[1] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs1_a2[2]$_SDFF_PN0_  (.D(_01033_),
    .Q(\CPU_rf_rd_index1_a2[2] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs1_a2[3]$_SDFF_PN0_  (.D(_01034_),
    .Q(\CPU_rf_rd_index1_a2[3] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs2_a2[0]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[20] ),
    .Q(\CPU_rf_rd_index2_a2[0] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs2_a2[1]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[21] ),
    .Q(\CPU_rf_rd_index2_a2[1] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs2_a2[2]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[22] ),
    .Q(\CPU_rf_rd_index2_a2[2] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_rs2_a2[3]$_DFF_P_  (.D(\CPU_imem_rd_data_a1[23] ),
    .Q(\CPU_rf_rd_index2_a2[3] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[0]$_DFF_P_  (.D(\CPU_src1_value_a2[0] ),
    .Q(\CPU_src1_value_a3[0] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src1_value_a3[10]$_DFF_P_  (.D(\CPU_src1_value_a2[10] ),
    .Q(\CPU_src1_value_a3[10] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src1_value_a3[11]$_DFF_P_  (.D(\CPU_src1_value_a2[11] ),
    .Q(\CPU_src1_value_a3[11] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[12]$_DFF_P_  (.D(\CPU_src1_value_a2[12] ),
    .Q(\CPU_src1_value_a3[12] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[13]$_DFF_P_  (.D(\CPU_src1_value_a2[13] ),
    .Q(\CPU_src1_value_a3[13] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[14]$_DFF_P_  (.D(\CPU_src1_value_a2[14] ),
    .Q(\CPU_src1_value_a3[14] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[15]$_DFF_P_  (.D(\CPU_src1_value_a2[15] ),
    .Q(\CPU_src1_value_a3[15] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[16]$_DFF_P_  (.D(\CPU_src1_value_a2[16] ),
    .Q(\CPU_src1_value_a3[16] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[17]$_DFF_P_  (.D(\CPU_src1_value_a2[17] ),
    .Q(\CPU_src1_value_a3[17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src1_value_a3[18]$_DFF_P_  (.D(\CPU_src1_value_a2[18] ),
    .Q(\CPU_src1_value_a3[18] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[19]$_DFF_P_  (.D(\CPU_src1_value_a2[19] ),
    .Q(\CPU_src1_value_a3[19] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[1]$_DFF_P_  (.D(\CPU_src1_value_a2[1] ),
    .Q(\CPU_src1_value_a3[1] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[20]$_DFF_P_  (.D(\CPU_src1_value_a2[20] ),
    .Q(\CPU_src1_value_a3[20] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[21]$_DFF_P_  (.D(\CPU_src1_value_a2[21] ),
    .Q(\CPU_src1_value_a3[21] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src1_value_a3[22]$_DFF_P_  (.D(\CPU_src1_value_a2[22] ),
    .Q(\CPU_src1_value_a3[22] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[23]$_DFF_P_  (.D(\CPU_src1_value_a2[23] ),
    .Q(\CPU_src1_value_a3[23] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[24]$_DFF_P_  (.D(\CPU_src1_value_a2[24] ),
    .Q(\CPU_src1_value_a3[24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[25]$_DFF_P_  (.D(\CPU_src1_value_a2[25] ),
    .Q(\CPU_src1_value_a3[25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[26]$_DFF_P_  (.D(\CPU_src1_value_a2[26] ),
    .Q(\CPU_src1_value_a3[26] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[27]$_DFF_P_  (.D(\CPU_src1_value_a2[27] ),
    .Q(\CPU_src1_value_a3[27] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[28]$_DFF_P_  (.D(\CPU_src1_value_a2[28] ),
    .Q(\CPU_src1_value_a3[28] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[29]$_DFF_P_  (.D(\CPU_src1_value_a2[29] ),
    .Q(\CPU_src1_value_a3[29] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[2]$_DFF_P_  (.D(\CPU_src1_value_a2[2] ),
    .Q(\CPU_src1_value_a3[2] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[30]$_DFF_P_  (.D(\CPU_src1_value_a2[30] ),
    .Q(\CPU_src1_value_a3[30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[31]$_DFF_P_  (.D(\CPU_src1_value_a2[31] ),
    .Q(\CPU_src1_value_a3[31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[3]$_DFF_P_  (.D(\CPU_src1_value_a2[3] ),
    .Q(\CPU_src1_value_a3[3] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[4]$_DFF_P_  (.D(\CPU_src1_value_a2[4] ),
    .Q(\CPU_src1_value_a3[4] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[5]$_DFF_P_  (.D(\CPU_src1_value_a2[5] ),
    .Q(\CPU_src1_value_a3[5] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[6]$_DFF_P_  (.D(\CPU_src1_value_a2[6] ),
    .Q(\CPU_src1_value_a3[6] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[7]$_DFF_P_  (.D(\CPU_src1_value_a2[7] ),
    .Q(\CPU_src1_value_a3[7] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src1_value_a3[8]$_DFF_P_  (.D(\CPU_src1_value_a2[8] ),
    .Q(\CPU_src1_value_a3[8] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src1_value_a3[9]$_DFF_P_  (.D(\CPU_src1_value_a2[9] ),
    .Q(\CPU_src1_value_a3[9] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[0]$_DFF_P_  (.D(\CPU_src2_value_a2[0] ),
    .Q(\CPU_src2_value_a3[0] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[10]$_DFF_P_  (.D(\CPU_src2_value_a2[10] ),
    .Q(\CPU_src2_value_a3[10] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[11]$_DFF_P_  (.D(\CPU_src2_value_a2[11] ),
    .Q(\CPU_src2_value_a3[11] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[12]$_DFF_P_  (.D(\CPU_src2_value_a2[12] ),
    .Q(\CPU_src2_value_a3[12] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a3[13]$_DFF_P_  (.D(\CPU_src2_value_a2[13] ),
    .Q(\CPU_src2_value_a3[13] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[14]$_DFF_P_  (.D(\CPU_src2_value_a2[14] ),
    .Q(\CPU_src2_value_a3[14] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[15]$_DFF_P_  (.D(\CPU_src2_value_a2[15] ),
    .Q(\CPU_src2_value_a3[15] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[16]$_DFF_P_  (.D(\CPU_src2_value_a2[16] ),
    .Q(\CPU_src2_value_a3[16] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[17]$_DFF_P_  (.D(\CPU_src2_value_a2[17] ),
    .Q(\CPU_src2_value_a3[17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[18]$_DFF_P_  (.D(\CPU_src2_value_a2[18] ),
    .Q(\CPU_src2_value_a3[18] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a3[19]$_DFF_P_  (.D(\CPU_src2_value_a2[19] ),
    .Q(\CPU_src2_value_a3[19] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[1]$_DFF_P_  (.D(\CPU_src2_value_a2[1] ),
    .Q(\CPU_src2_value_a3[1] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[20]$_DFF_P_  (.D(\CPU_src2_value_a2[20] ),
    .Q(\CPU_src2_value_a3[20] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[21]$_DFF_P_  (.D(\CPU_src2_value_a2[21] ),
    .Q(\CPU_src2_value_a3[21] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[22]$_DFF_P_  (.D(\CPU_src2_value_a2[22] ),
    .Q(\CPU_src2_value_a3[22] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a3[23]$_DFF_P_  (.D(\CPU_src2_value_a2[23] ),
    .Q(\CPU_src2_value_a3[23] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[24]$_DFF_P_  (.D(\CPU_src2_value_a2[24] ),
    .Q(\CPU_src2_value_a3[24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[25]$_DFF_P_  (.D(\CPU_src2_value_a2[25] ),
    .Q(\CPU_src2_value_a3[25] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[26]$_DFF_P_  (.D(\CPU_src2_value_a2[26] ),
    .Q(\CPU_src2_value_a3[26] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[27]$_DFF_P_  (.D(\CPU_src2_value_a2[27] ),
    .Q(\CPU_src2_value_a3[27] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[28]$_DFF_P_  (.D(\CPU_src2_value_a2[28] ),
    .Q(\CPU_src2_value_a3[28] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[29]$_DFF_P_  (.D(\CPU_src2_value_a2[29] ),
    .Q(\CPU_src2_value_a3[29] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[2]$_DFF_P_  (.D(\CPU_src2_value_a2[2] ),
    .Q(\CPU_src2_value_a3[2] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[30]$_DFF_P_  (.D(\CPU_src2_value_a2[30] ),
    .Q(\CPU_src2_value_a3[30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[31]$_DFF_P_  (.D(\CPU_src2_value_a2[31] ),
    .Q(\CPU_src2_value_a3[31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[3]$_DFF_P_  (.D(\CPU_src2_value_a2[3] ),
    .Q(\CPU_src2_value_a3[3] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[4]$_DFF_P_  (.D(\CPU_src2_value_a2[4] ),
    .Q(\CPU_src2_value_a3[4] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[5]$_DFF_P_  (.D(\CPU_src2_value_a2[5] ),
    .Q(\CPU_src2_value_a3[5] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[6]$_DFF_P_  (.D(\CPU_src2_value_a2[6] ),
    .Q(\CPU_src2_value_a3[6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_src2_value_a3[7]$_DFF_P_  (.D(\CPU_src2_value_a2[7] ),
    .Q(\CPU_src2_value_a3[7] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[8]$_DFF_P_  (.D(\CPU_src2_value_a2[8] ),
    .Q(\CPU_src2_value_a3[8] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 \CPU_src2_value_a3[9]$_DFF_P_  (.D(\CPU_src2_value_a2[9] ),
    .Q(\CPU_src2_value_a3[9] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[0]$_DFF_P_  (.D(net184),
    .Q(\CPU_dmem_wr_data_a4[0] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[10]$_DFF_P_  (.D(net176),
    .Q(\CPU_dmem_wr_data_a4[10] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[11]$_DFF_P_  (.D(net190),
    .Q(\CPU_dmem_wr_data_a4[11] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[12]$_DFF_P_  (.D(net181),
    .Q(\CPU_dmem_wr_data_a4[12] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[13]$_DFF_P_  (.D(net702),
    .Q(\CPU_dmem_wr_data_a4[13] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[14]$_DFF_P_  (.D(net178),
    .Q(\CPU_dmem_wr_data_a4[14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[15]$_DFF_P_  (.D(net599),
    .Q(\CPU_dmem_wr_data_a4[15] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[16]$_DFF_P_  (.D(net198),
    .Q(\CPU_dmem_wr_data_a4[16] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[17]$_DFF_P_  (.D(net185),
    .Q(\CPU_dmem_wr_data_a4[17] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[18]$_DFF_P_  (.D(net201),
    .Q(\CPU_dmem_wr_data_a4[18] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[19]$_DFF_P_  (.D(net194),
    .Q(\CPU_dmem_wr_data_a4[19] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[1]$_DFF_P_  (.D(net164),
    .Q(\CPU_dmem_wr_data_a4[1] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[20]$_DFF_P_  (.D(net199),
    .Q(\CPU_dmem_wr_data_a4[20] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[21]$_DFF_P_  (.D(net200),
    .Q(\CPU_dmem_wr_data_a4[21] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[22]$_DFF_P_  (.D(net183),
    .Q(\CPU_dmem_wr_data_a4[22] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[23]$_DFF_P_  (.D(net214),
    .Q(\CPU_dmem_wr_data_a4[23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[24]$_DFF_P_  (.D(net162),
    .Q(\CPU_dmem_wr_data_a4[24] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[25]$_DFF_P_  (.D(net173),
    .Q(\CPU_dmem_wr_data_a4[25] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[26]$_DFF_P_  (.D(net163),
    .Q(\CPU_dmem_wr_data_a4[26] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[27]$_DFF_P_  (.D(net193),
    .Q(\CPU_dmem_wr_data_a4[27] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[28]$_DFF_P_  (.D(net196),
    .Q(\CPU_dmem_wr_data_a4[28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[29]$_DFF_P_  (.D(net175),
    .Q(\CPU_dmem_wr_data_a4[29] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[2]$_DFF_P_  (.D(net169),
    .Q(\CPU_dmem_wr_data_a4[2] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[30]$_DFF_P_  (.D(net167),
    .Q(\CPU_dmem_wr_data_a4[30] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[31]$_DFF_P_  (.D(net917),
    .Q(\CPU_dmem_wr_data_a4[31] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[3]$_DFF_P_  (.D(net160),
    .Q(\CPU_dmem_wr_data_a4[3] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[4]$_DFF_P_  (.D(net170),
    .Q(\CPU_dmem_wr_data_a4[4] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[5]$_DFF_P_  (.D(net188),
    .Q(\CPU_dmem_wr_data_a4[5] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[6]$_DFF_P_  (.D(net197),
    .Q(\CPU_dmem_wr_data_a4[6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[7]$_DFF_P_  (.D(net189),
    .Q(\CPU_dmem_wr_data_a4[7] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[8]$_DFF_P_  (.D(net439),
    .Q(\CPU_dmem_wr_data_a4[8] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_4 \CPU_src2_value_a4[9]$_DFF_P_  (.D(net187),
    .Q(\CPU_dmem_wr_data_a4[9] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_valid_a4$_DFF_P_  (.D(_01036_),
    .Q(CPU_valid_a4),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_valid_load_a4$_DFF_P_  (.D(CPU_valid_load_a3),
    .Q(CPU_dmem_rd_en_a4),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_valid_load_a5$_DFF_P_  (.D(net151),
    .Q(CPU_valid_load_a5),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_valid_taken_br_a4$_DFF_P_  (.D(CPU_valid_taken_br_a3),
    .Q(CPU_valid_taken_br_a4),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 \CPU_valid_taken_br_a5$_DFF_P_  (.D(net147),
    .Q(CPU_valid_taken_br_a5),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__or4_4 _05825_ (.A(CPU_valid_load_a5),
    .B(CPU_valid_taken_br_a5),
    .C(CPU_valid_taken_br_a4),
    .D(CPU_dmem_rd_en_a4),
    .X(_01035_));
 sky130_fd_sc_hd__clkinv_16 _05826_ (.A(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_672 ();
 sky130_fd_sc_hd__a21o_1 _05831_ (.A1(_05790_),
    .A2(_05795_),
    .B1(_05794_),
    .X(_01040_));
 sky130_fd_sc_hd__a21o_1 _05832_ (.A1(_05804_),
    .A2(_01040_),
    .B1(_05803_),
    .X(_01041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_671 ();
 sky130_fd_sc_hd__nand4_2 _05834_ (.A(_05525_),
    .B(_05791_),
    .C(_05795_),
    .D(_05804_),
    .Y(_01043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_669 ();
 sky130_fd_sc_hd__inv_1 _05837_ (.A(_05787_),
    .Y(_01046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_668 ();
 sky130_fd_sc_hd__a21oi_1 _05839_ (.A1(_05773_),
    .A2(_05778_),
    .B1(_05777_),
    .Y(_01048_));
 sky130_fd_sc_hd__o21bai_1 _05840_ (.A1(_01046_),
    .A2(_01048_),
    .B1_N(_05786_),
    .Y(_01049_));
 sky130_fd_sc_hd__a21oi_2 _05841_ (.A1(_05528_),
    .A2(_01049_),
    .B1(_05527_),
    .Y(_01050_));
 sky130_fd_sc_hd__nor2_1 _05842_ (.A(_01043_),
    .B(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__a211oi_4 _05843_ (.A1(_05525_),
    .A2(_01041_),
    .B1(_01051_),
    .C1(_05524_),
    .Y(_01052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_667 ();
 sky130_fd_sc_hd__nand4_1 _05845_ (.A(_05543_),
    .B(_05708_),
    .C(_05717_),
    .D(_05726_),
    .Y(_01054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_664 ();
 sky130_fd_sc_hd__a21o_1 _05849_ (.A1(_05680_),
    .A2(_05690_),
    .B1(_05689_),
    .X(_01058_));
 sky130_fd_sc_hd__a21o_1 _05850_ (.A1(_05699_),
    .A2(_01058_),
    .B1(_05698_),
    .X(_01059_));
 sky130_fd_sc_hd__a21oi_1 _05851_ (.A1(_05548_),
    .A2(_01059_),
    .B1(_05547_),
    .Y(_01060_));
 sky130_fd_sc_hd__inv_1 _05852_ (.A(_05726_),
    .Y(_01061_));
 sky130_fd_sc_hd__a21oi_1 _05853_ (.A1(_05707_),
    .A2(_05717_),
    .B1(_05716_),
    .Y(_01062_));
 sky130_fd_sc_hd__o21bai_1 _05854_ (.A1(_01061_),
    .A2(_01062_),
    .B1_N(_05725_),
    .Y(_01063_));
 sky130_fd_sc_hd__a21oi_1 _05855_ (.A1(_05543_),
    .A2(_01063_),
    .B1(_05542_),
    .Y(_01064_));
 sky130_fd_sc_hd__inv_1 _05856_ (.A(_05538_),
    .Y(_01065_));
 sky130_fd_sc_hd__inv_1 _05857_ (.A(_05752_),
    .Y(_01066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_662 ();
 sky130_fd_sc_hd__a21o_1 _05860_ (.A1(_05729_),
    .A2(_05734_),
    .B1(_05733_),
    .X(_01069_));
 sky130_fd_sc_hd__a21oi_1 _05861_ (.A1(_05743_),
    .A2(_01069_),
    .B1(_05742_),
    .Y(_01070_));
 sky130_fd_sc_hd__a21oi_1 _05862_ (.A1(_05752_),
    .A2(_05537_),
    .B1(_05751_),
    .Y(_01071_));
 sky130_fd_sc_hd__o31a_1 _05863_ (.A1(_01065_),
    .A2(_01066_),
    .A3(_01070_),
    .B1(_01071_),
    .X(_01072_));
 sky130_fd_sc_hd__o211ai_1 _05864_ (.A1(_01054_),
    .A2(_01060_),
    .B1(_01064_),
    .C1(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__and3_1 _05865_ (.A(_05538_),
    .B(_05730_),
    .C(_05734_),
    .X(_01074_));
 sky130_fd_sc_hd__nand3_1 _05866_ (.A(_05743_),
    .B(_05752_),
    .C(_01074_),
    .Y(_01075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_660 ();
 sky130_fd_sc_hd__nand3_2 _05869_ (.A(_05533_),
    .B(_05761_),
    .C(_05770_),
    .Y(_01078_));
 sky130_fd_sc_hd__a21oi_1 _05870_ (.A1(_01072_),
    .A2(_01075_),
    .B1(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hd__clkinvlp_4 _05871_ (.A(_05553_),
    .Y(_01080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_659 ();
 sky130_fd_sc_hd__nor2_1 _05873_ (.A(_05672_),
    .B(_05671_),
    .Y(_01082_));
 sky130_fd_sc_hd__nor2_1 _05874_ (.A(_01080_),
    .B(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__nor2_1 _05875_ (.A(_05552_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_657 ();
 sky130_fd_sc_hd__nand4_1 _05878_ (.A(_05558_),
    .B(_05645_),
    .C(_05654_),
    .D(_05663_),
    .Y(_01087_));
 sky130_fd_sc_hd__inv_1 _05879_ (.A(_05635_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21oi_1 _05880_ (.A1(_05562_),
    .A2(_01088_),
    .B1(_05561_),
    .Y(_01089_));
 sky130_fd_sc_hd__a21o_1 _05881_ (.A1(_05558_),
    .A2(_05644_),
    .B1(_05557_),
    .X(_01090_));
 sky130_fd_sc_hd__nand3_1 _05882_ (.A(_05654_),
    .B(_05663_),
    .C(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__a211oi_1 _05883_ (.A1(_05553_),
    .A2(_05671_),
    .B1(_05662_),
    .C1(_05552_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _05884_ (.A(_05653_),
    .B(_05663_),
    .Y(_01093_));
 sky130_fd_sc_hd__o2111a_1 _05885_ (.A1(_01087_),
    .A2(_01089_),
    .B1(_01091_),
    .C1(_01092_),
    .D1(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__nand4_1 _05886_ (.A(_05548_),
    .B(_05681_),
    .C(_05690_),
    .D(_05699_),
    .Y(_01095_));
 sky130_fd_sc_hd__or4_1 _05887_ (.A(_01078_),
    .B(_01075_),
    .C(_01054_),
    .D(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__inv_1 _05888_ (.A(_05533_),
    .Y(_01097_));
 sky130_fd_sc_hd__a21oi_1 _05889_ (.A1(_05770_),
    .A2(_05760_),
    .B1(_05769_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _05890_ (.A(_01097_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _05891_ (.A(_05532_),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__o31ai_1 _05892_ (.A1(_01084_),
    .A2(_01094_),
    .A3(_01096_),
    .B1(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__a21oi_1 _05893_ (.A1(_01073_),
    .A2(_01079_),
    .B1(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand4_1 _05894_ (.A(_05528_),
    .B(_05774_),
    .C(_05778_),
    .D(_05787_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_2 _05895_ (.A(_01043_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__a211oi_1 _05896_ (.A1(_05525_),
    .A2(_01041_),
    .B1(_01104_),
    .C1(_05524_),
    .Y(_01105_));
 sky130_fd_sc_hd__o21ai_2 _05897_ (.A1(_01043_),
    .A2(_01050_),
    .B1(_01105_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand4_1 _05898_ (.A(_05553_),
    .B(_05562_),
    .C(_05636_),
    .D(_05672_),
    .Y(_01107_));
 sky130_fd_sc_hd__nor2_1 _05899_ (.A(_01087_),
    .B(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3b_1 _05900_ (.A_N(_01096_),
    .B(_01104_),
    .C(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _05901_ (.A(_01106_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__a21oi_1 _05902_ (.A1(_01052_),
    .A2(_01102_),
    .B1(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__nand2_1 _05903_ (.A(_05525_),
    .B(CPU_is_blt_a3),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2b_1 _05904_ (.A_N(CPU_is_blt_a3),
    .B(CPU_is_bltu_a3),
    .Y(_01113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_655 ();
 sky130_fd_sc_hd__a21oi_1 _05907_ (.A1(_01112_),
    .A2(_01113_),
    .B1(_01035_),
    .Y(_01116_));
 sky130_fd_sc_hd__and4b_1 _05908_ (.A_N(_05525_),
    .B(CPU_is_blt_a3),
    .C(_01036_),
    .D(_01110_),
    .X(_01117_));
 sky130_fd_sc_hd__a21oi_4 _05909_ (.A1(_01111_),
    .A2(_01116_),
    .B1(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__inv_1 _05910_ (.A(_01118_),
    .Y(CPU_valid_taken_br_a3));
 sky130_fd_sc_hd__nand2_4 _05911_ (.A(net1831),
    .B(_01036_),
    .Y(_01119_));
 sky130_fd_sc_hd__inv_1 _05912_ (.A(_01119_),
    .Y(CPU_valid_load_a3));
 sky130_fd_sc_hd__inv_1 _05913_ (.A(net1569),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_1 _05914_ (.A(_01120_),
    .B(net1833),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _05915_ (.A(_05818_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__inv_1 _05916_ (.A(_01122_),
    .Y(\CPU_dec_bits_a1[10] ));
 sky130_fd_sc_hd__inv_1 _05917_ (.A(net192),
    .Y(\CPU_inc_pc_a1[2] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_653 ();
 sky130_fd_sc_hd__xor2_1 _05920_ (.A(net827),
    .B(_05822_),
    .X(\CPU_inc_pc_a1[4] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_652 ();
 sky130_fd_sc_hd__nand3_1 _05922_ (.A(net827),
    .B(net182),
    .C(net192),
    .Y(_01126_));
 sky130_fd_sc_hd__xnor2_1 _05923_ (.A(net1291),
    .B(_01126_),
    .Y(\CPU_inc_pc_a1[5] ));
 sky130_fd_sc_hd__a21oi_1 _05924_ (.A1(\CPU_imem_rd_addr_a1[3] ),
    .A2(_05817_),
    .B1(_05820_),
    .Y(_01127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_651 ();
 sky130_fd_sc_hd__inv_1 _05926_ (.A(_05820_),
    .Y(_01129_));
 sky130_fd_sc_hd__nor2_1 _05927_ (.A(_05818_),
    .B(_05822_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _05928_ (.A(_01129_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__a21oi_1 _05929_ (.A1(net827),
    .A2(_05817_),
    .B1(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__o32ai_2 _05930_ (.A1(net1569),
    .A2(net182),
    .A3(_01127_),
    .B1(_01132_),
    .B2(net1833),
    .Y(_01133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_650 ();
 sky130_fd_sc_hd__nor3_1 _05932_ (.A(\CPU_imem_rd_addr_a1[2] ),
    .B(\CPU_imem_rd_addr_a1[3] ),
    .C(_05822_),
    .Y(_01135_));
 sky130_fd_sc_hd__a21oi_1 _05933_ (.A1(net1847),
    .A2(_01129_),
    .B1(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_649 ();
 sky130_fd_sc_hd__nor2_1 _05935_ (.A(_05818_),
    .B(_05820_),
    .Y(_01138_));
 sky130_fd_sc_hd__o21ai_0 _05936_ (.A1(net1847),
    .A2(_01138_),
    .B1(net827),
    .Y(_01139_));
 sky130_fd_sc_hd__nand3_1 _05937_ (.A(_01133_),
    .B(_01136_),
    .C(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__inv_1 _05938_ (.A(_01140_),
    .Y(\CPU_imem_rd_data_a1[7] ));
 sky130_fd_sc_hd__inv_1 _05939_ (.A(_05817_),
    .Y(_01141_));
 sky130_fd_sc_hd__a21oi_1 _05940_ (.A1(_01141_),
    .A2(_05820_),
    .B1(\CPU_imem_rd_addr_a1[1] ),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_1 _05941_ (.A(_05822_),
    .B(_05820_),
    .Y(_01143_));
 sky130_fd_sc_hd__a21oi_1 _05942_ (.A1(_05818_),
    .A2(_01143_),
    .B1(\CPU_imem_rd_addr_a1[3] ),
    .Y(_01144_));
 sky130_fd_sc_hd__a21oi_1 _05943_ (.A1(\CPU_imem_rd_addr_a1[3] ),
    .A2(_01142_),
    .B1(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__and3_1 _05944_ (.A(_01141_),
    .B(_05820_),
    .C(_01130_),
    .X(_01146_));
 sky130_fd_sc_hd__nand2b_1 _05945_ (.A_N(net1833),
    .B(net827),
    .Y(_01147_));
 sky130_fd_sc_hd__o22a_1 _05946_ (.A1(net1851),
    .A2(_01145_),
    .B1(_01146_),
    .B2(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__nor4_1 _05947_ (.A(_05822_),
    .B(_05817_),
    .C(_05820_),
    .D(_01122_),
    .Y(\CPU_imm_a1[10] ));
 sky130_fd_sc_hd__nor2_1 _05948_ (.A(_05817_),
    .B(_05820_),
    .Y(_01149_));
 sky130_fd_sc_hd__nor3b_1 _05949_ (.A(net1569),
    .B(_01149_),
    .C_N(\CPU_imem_rd_addr_a1[3] ),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _05950_ (.A(\CPU_imm_a1[10] ),
    .B(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _05951_ (.A(_01148_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _05952_ (.A(_01122_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__inv_1 _05953_ (.A(_01153_),
    .Y(CPU_is_s_instr_a1));
 sky130_fd_sc_hd__or4_1 _05954_ (.A(_01120_),
    .B(_05822_),
    .C(_05817_),
    .D(_01138_),
    .X(_01154_));
 sky130_fd_sc_hd__o31ai_1 _05955_ (.A1(net827),
    .A2(_05820_),
    .A3(_01130_),
    .B1(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _05956_ (.A(net1569),
    .B(net182),
    .Y(_01156_));
 sky130_fd_sc_hd__o21ai_1 _05957_ (.A1(_01141_),
    .A2(_05820_),
    .B1(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__mux2i_1 _05958_ (.A0(_01155_),
    .A1(_01157_),
    .S(net1291),
    .Y(\CPU_imem_rd_data_a1[8] ));
 sky130_fd_sc_hd__o21ai_0 _05959_ (.A1(net182),
    .A2(_01149_),
    .B1(net1291),
    .Y(_01158_));
 sky130_fd_sc_hd__o21ai_0 _05960_ (.A1(net1833),
    .A2(_01149_),
    .B1(net827),
    .Y(_01159_));
 sky130_fd_sc_hd__o311a_1 _05961_ (.A1(net827),
    .A2(net1291),
    .A3(_01131_),
    .B1(_01158_),
    .C1(_01159_),
    .X(\CPU_imem_rd_data_a1[9] ));
 sky130_fd_sc_hd__nand2_1 _05962_ (.A(net1291),
    .B(_01157_),
    .Y(\CPU_imem_rd_data_a1[10] ));
 sky130_fd_sc_hd__inv_1 _05963_ (.A(\CPU_imm_a3[1] ),
    .Y(_05510_));
 sky130_fd_sc_hd__inv_1 _05964_ (.A(net159),
    .Y(_05519_));
 sky130_fd_sc_hd__inv_1 _05965_ (.A(\CPU_src2_value_a3[1] ),
    .Y(_05515_));
 sky130_fd_sc_hd__inv_1 _05966_ (.A(net156),
    .Y(_05520_));
 sky130_fd_sc_hd__inv_1 _05967_ (.A(_05630_),
    .Y(_05512_));
 sky130_fd_sc_hd__inv_1 _05968_ (.A(_05637_),
    .Y(_05516_));
 sky130_fd_sc_hd__inv_1 _05969_ (.A(_05815_),
    .Y(_05521_));
 sky130_fd_sc_hd__inv_1 _05970_ (.A(\CPU_imm_a3[0] ),
    .Y(_05627_));
 sky130_fd_sc_hd__inv_1 _05971_ (.A(\CPU_src1_value_a3[2] ),
    .Y(_05639_));
 sky130_fd_sc_hd__inv_1 _05972_ (.A(\CPU_src1_value_a3[4] ),
    .Y(_05648_));
 sky130_fd_sc_hd__inv_1 _05973_ (.A(\CPU_src1_value_a3[5] ),
    .Y(_05657_));
 sky130_fd_sc_hd__inv_1 _05974_ (.A(\CPU_src1_value_a3[6] ),
    .Y(_05666_));
 sky130_fd_sc_hd__inv_1 _05975_ (.A(\CPU_src1_value_a3[8] ),
    .Y(_05675_));
 sky130_fd_sc_hd__inv_1 _05976_ (.A(\CPU_src1_value_a3[9] ),
    .Y(_05684_));
 sky130_fd_sc_hd__inv_1 _05977_ (.A(\CPU_src1_value_a3[10] ),
    .Y(_05693_));
 sky130_fd_sc_hd__inv_1 _05978_ (.A(\CPU_src1_value_a3[12] ),
    .Y(_05702_));
 sky130_fd_sc_hd__inv_1 _05979_ (.A(\CPU_src1_value_a3[13] ),
    .Y(_05711_));
 sky130_fd_sc_hd__inv_1 _05980_ (.A(\CPU_src1_value_a3[14] ),
    .Y(_05720_));
 sky130_fd_sc_hd__inv_1 _05981_ (.A(\CPU_src1_value_a3[16] ),
    .Y(_05602_));
 sky130_fd_sc_hd__inv_1 _05982_ (.A(\CPU_src1_value_a3[17] ),
    .Y(_05597_));
 sky130_fd_sc_hd__inv_1 _05983_ (.A(\CPU_src1_value_a3[18] ),
    .Y(_05737_));
 sky130_fd_sc_hd__inv_1 _05984_ (.A(\CPU_src1_value_a3[20] ),
    .Y(_05746_));
 sky130_fd_sc_hd__inv_1 _05985_ (.A(\CPU_src1_value_a3[21] ),
    .Y(_05755_));
 sky130_fd_sc_hd__inv_1 _05986_ (.A(\CPU_src1_value_a3[22] ),
    .Y(_05764_));
 sky130_fd_sc_hd__inv_1 _05987_ (.A(\CPU_src1_value_a3[24] ),
    .Y(_05584_));
 sky130_fd_sc_hd__inv_1 _05988_ (.A(\CPU_src1_value_a3[25] ),
    .Y(_05579_));
 sky130_fd_sc_hd__inv_1 _05989_ (.A(\CPU_src1_value_a3[26] ),
    .Y(_05781_));
 sky130_fd_sc_hd__inv_1 _05990_ (.A(\CPU_src1_value_a3[28] ),
    .Y(_05570_));
 sky130_fd_sc_hd__inv_1 _05991_ (.A(\CPU_src1_value_a3[29] ),
    .Y(_05565_));
 sky130_fd_sc_hd__inv_1 _05992_ (.A(\CPU_src1_value_a3[30] ),
    .Y(_05798_));
 sky130_fd_sc_hd__inv_1 _05993_ (.A(\CPU_src1_value_a3[27] ),
    .Y(_05526_));
 sky130_fd_sc_hd__inv_1 _05994_ (.A(\CPU_src1_value_a3[23] ),
    .Y(_05531_));
 sky130_fd_sc_hd__inv_1 _05995_ (.A(\CPU_src1_value_a3[19] ),
    .Y(_05536_));
 sky130_fd_sc_hd__inv_1 _05996_ (.A(\CPU_src1_value_a3[15] ),
    .Y(_05541_));
 sky130_fd_sc_hd__inv_1 _05997_ (.A(\CPU_src1_value_a3[11] ),
    .Y(_05546_));
 sky130_fd_sc_hd__inv_1 _05998_ (.A(\CPU_src1_value_a3[7] ),
    .Y(_05551_));
 sky130_fd_sc_hd__inv_1 _05999_ (.A(\CPU_src1_value_a3[3] ),
    .Y(_05556_));
 sky130_fd_sc_hd__clkinvlp_4 _06000_ (.A(\CPU_src1_value_a3[1] ),
    .Y(_05511_));
 sky130_fd_sc_hd__clkinv_4 _06001_ (.A(\CPU_src1_value_a3[31] ),
    .Y(_05523_));
 sky130_fd_sc_hd__inv_1 _06002_ (.A(\CPU_src2_value_a3[0] ),
    .Y(_05634_));
 sky130_fd_sc_hd__inv_1 _06003_ (.A(net182),
    .Y(_05816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_647 ();
 sky130_fd_sc_hd__nand2_8 _06006_ (.A(CPU_is_s_instr_a4),
    .B(CPU_valid_a4),
    .Y(_01162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_644 ();
 sky130_fd_sc_hd__nor2_2 _06010_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .Y(_01166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_642 ();
 sky130_fd_sc_hd__nor2_2 _06013_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_8 _06014_ (.A(_01166_),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__nor2_8 _06015_ (.A(_01162_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_641 ();
 sky130_fd_sc_hd__nand2_1 _06017_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(_01171_),
    .Y(_01173_));
 sky130_fd_sc_hd__and2_4 _06018_ (.A(CPU_is_s_instr_a4),
    .B(CPU_valid_a4),
    .X(_01174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_639 ();
 sky130_fd_sc_hd__nor4_4 _06021_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(\CPU_dmem_addr_a4[2] ),
    .D(\CPU_dmem_addr_a4[3] ),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_8 _06022_ (.A(_01174_),
    .B(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_638 ();
 sky130_fd_sc_hd__nand2_1 _06024_ (.A(net848),
    .B(_01178_),
    .Y(_01180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_635 ();
 sky130_fd_sc_hd__a21oi_1 _06028_ (.A1(_01173_),
    .A2(_01180_),
    .B1(net104),
    .Y(_00000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_633 ();
 sky130_fd_sc_hd__nand2_1 _06031_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(_01171_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _06032_ (.A(net500),
    .B(_01178_),
    .Y(_01187_));
 sky130_fd_sc_hd__a21oi_1 _06033_ (.A1(_01186_),
    .A2(_01187_),
    .B1(net107),
    .Y(_00001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_631 ();
 sky130_fd_sc_hd__nand2_1 _06036_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(_01171_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _06037_ (.A(net299),
    .B(_01178_),
    .Y(_01191_));
 sky130_fd_sc_hd__a21oi_1 _06038_ (.A1(_01190_),
    .A2(_01191_),
    .B1(net106),
    .Y(_00002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_629 ();
 sky130_fd_sc_hd__nand2_1 _06041_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(_01171_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _06042_ (.A(net371),
    .B(_01178_),
    .Y(_01195_));
 sky130_fd_sc_hd__a21oi_1 _06043_ (.A1(_01194_),
    .A2(_01195_),
    .B1(net107),
    .Y(_00003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_627 ();
 sky130_fd_sc_hd__nand2_1 _06046_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(_01171_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _06047_ (.A(net537),
    .B(_01178_),
    .Y(_01199_));
 sky130_fd_sc_hd__a21oi_1 _06048_ (.A1(_01198_),
    .A2(_01199_),
    .B1(net106),
    .Y(_00004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_625 ();
 sky130_fd_sc_hd__nand2_1 _06051_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(_01171_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _06052_ (.A(net315),
    .B(_01178_),
    .Y(_01203_));
 sky130_fd_sc_hd__a21oi_1 _06053_ (.A1(_01202_),
    .A2(_01203_),
    .B1(net107),
    .Y(_00005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_623 ();
 sky130_fd_sc_hd__nand2_1 _06056_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(_01171_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _06057_ (.A(net472),
    .B(_01178_),
    .Y(_01207_));
 sky130_fd_sc_hd__a21oi_1 _06058_ (.A1(_01206_),
    .A2(_01207_),
    .B1(net104),
    .Y(_00006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_621 ();
 sky130_fd_sc_hd__nand2_1 _06061_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(_01171_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _06062_ (.A(net1162),
    .B(_01178_),
    .Y(_01211_));
 sky130_fd_sc_hd__a21oi_1 _06063_ (.A1(_01210_),
    .A2(_01211_),
    .B1(net105),
    .Y(_00007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_619 ();
 sky130_fd_sc_hd__nand2_1 _06066_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(_01171_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_1 _06067_ (.A(net741),
    .B(_01178_),
    .Y(_01215_));
 sky130_fd_sc_hd__a21oi_1 _06068_ (.A1(_01214_),
    .A2(_01215_),
    .B1(net102),
    .Y(_00008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_617 ();
 sky130_fd_sc_hd__nand2_1 _06071_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(_01171_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand2_1 _06072_ (.A(net1018),
    .B(_01178_),
    .Y(_01219_));
 sky130_fd_sc_hd__a21oi_1 _06073_ (.A1(_01218_),
    .A2(_01219_),
    .B1(net106),
    .Y(_00009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_614 ();
 sky130_fd_sc_hd__nand2_1 _06077_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(_01171_),
    .Y(_01223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_613 ();
 sky130_fd_sc_hd__nand2_1 _06079_ (.A(net543),
    .B(_01178_),
    .Y(_01225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_612 ();
 sky130_fd_sc_hd__a21oi_1 _06081_ (.A1(_01223_),
    .A2(_01225_),
    .B1(net106),
    .Y(_00010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_610 ();
 sky130_fd_sc_hd__nand2_1 _06084_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01171_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _06085_ (.A(net387),
    .B(_01178_),
    .Y(_01230_));
 sky130_fd_sc_hd__a21oi_1 _06086_ (.A1(_01229_),
    .A2(_01230_),
    .B1(net103),
    .Y(_00011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_608 ();
 sky130_fd_sc_hd__nand2_1 _06089_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(_01171_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _06090_ (.A(net646),
    .B(_01178_),
    .Y(_01234_));
 sky130_fd_sc_hd__a21oi_1 _06091_ (.A1(_01233_),
    .A2(_01234_),
    .B1(net102),
    .Y(_00012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_606 ();
 sky130_fd_sc_hd__nand2_1 _06094_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(_01171_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _06095_ (.A(net838),
    .B(_01178_),
    .Y(_01238_));
 sky130_fd_sc_hd__a21oi_1 _06096_ (.A1(_01237_),
    .A2(_01238_),
    .B1(net104),
    .Y(_00013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_604 ();
 sky130_fd_sc_hd__nand2_1 _06099_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(_01171_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _06100_ (.A(net1077),
    .B(_01178_),
    .Y(_01242_));
 sky130_fd_sc_hd__a21oi_1 _06101_ (.A1(_01241_),
    .A2(_01242_),
    .B1(net106),
    .Y(_00014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_602 ();
 sky130_fd_sc_hd__nand2_1 _06104_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_01171_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(net775),
    .B(_01178_),
    .Y(_01246_));
 sky130_fd_sc_hd__a21oi_1 _06106_ (.A1(_01245_),
    .A2(_01246_),
    .B1(net102),
    .Y(_00015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_600 ();
 sky130_fd_sc_hd__nand2_1 _06109_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(_01171_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _06110_ (.A(net383),
    .B(_01178_),
    .Y(_01250_));
 sky130_fd_sc_hd__a21oi_1 _06111_ (.A1(_01249_),
    .A2(_01250_),
    .B1(CPU_reset_a4),
    .Y(_00016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_598 ();
 sky130_fd_sc_hd__nand2_1 _06114_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(_01171_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _06115_ (.A(net553),
    .B(_01178_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21oi_1 _06116_ (.A1(_01253_),
    .A2(_01254_),
    .B1(net106),
    .Y(_00017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_596 ();
 sky130_fd_sc_hd__nand2_1 _06119_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(_01171_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(net1075),
    .B(_01178_),
    .Y(_01258_));
 sky130_fd_sc_hd__a21oi_1 _06121_ (.A1(_01257_),
    .A2(_01258_),
    .B1(net107),
    .Y(_00018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_594 ();
 sky130_fd_sc_hd__nand2_1 _06124_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(_01171_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2_1 _06125_ (.A(net844),
    .B(_01178_),
    .Y(_01262_));
 sky130_fd_sc_hd__a21oi_1 _06126_ (.A1(_01261_),
    .A2(_01262_),
    .B1(net105),
    .Y(_00019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_591 ();
 sky130_fd_sc_hd__nand2_1 _06130_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(_01171_),
    .Y(_01266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_590 ();
 sky130_fd_sc_hd__nand2_1 _06132_ (.A(net753),
    .B(_01178_),
    .Y(_01268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_589 ();
 sky130_fd_sc_hd__a21oi_1 _06134_ (.A1(_01266_),
    .A2(_01268_),
    .B1(net104),
    .Y(_00020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_587 ();
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(_01171_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _06138_ (.A(net369),
    .B(_01178_),
    .Y(_01273_));
 sky130_fd_sc_hd__a21oi_1 _06139_ (.A1(_01272_),
    .A2(_01273_),
    .B1(net107),
    .Y(_00021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_585 ();
 sky130_fd_sc_hd__nand2_1 _06142_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01171_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _06143_ (.A(net399),
    .B(_01178_),
    .Y(_01277_));
 sky130_fd_sc_hd__a21oi_1 _06144_ (.A1(_01276_),
    .A2(_01277_),
    .B1(net103),
    .Y(_00022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_583 ();
 sky130_fd_sc_hd__nand2_1 _06147_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(_01171_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _06148_ (.A(net1083),
    .B(_01178_),
    .Y(_01281_));
 sky130_fd_sc_hd__a21oi_1 _06149_ (.A1(_01280_),
    .A2(_01281_),
    .B1(net107),
    .Y(_00023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_581 ();
 sky130_fd_sc_hd__nand2_1 _06152_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(_01171_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _06153_ (.A(net450),
    .B(_01178_),
    .Y(_01285_));
 sky130_fd_sc_hd__a21oi_1 _06154_ (.A1(_01284_),
    .A2(_01285_),
    .B1(net105),
    .Y(_00024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_579 ();
 sky130_fd_sc_hd__nand2_1 _06157_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01171_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _06158_ (.A(net992),
    .B(_01178_),
    .Y(_01289_));
 sky130_fd_sc_hd__a21oi_1 _06159_ (.A1(_01288_),
    .A2(_01289_),
    .B1(net103),
    .Y(_00025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_577 ();
 sky130_fd_sc_hd__nand2_1 _06162_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_01171_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _06163_ (.A(net729),
    .B(_01178_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21oi_1 _06164_ (.A1(_01292_),
    .A2(_01293_),
    .B1(net103),
    .Y(_00026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_575 ();
 sky130_fd_sc_hd__nand2_1 _06167_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01171_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(net488),
    .B(_01178_),
    .Y(_01297_));
 sky130_fd_sc_hd__a21oi_1 _06169_ (.A1(_01296_),
    .A2(_01297_),
    .B1(net105),
    .Y(_00027_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_573 ();
 sky130_fd_sc_hd__nand2_1 _06172_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(_01171_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _06173_ (.A(net890),
    .B(_01178_),
    .Y(_01301_));
 sky130_fd_sc_hd__a21oi_1 _06174_ (.A1(_01300_),
    .A2(_01301_),
    .B1(net107),
    .Y(_00028_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_571 ();
 sky130_fd_sc_hd__nand2_1 _06177_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_01171_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _06178_ (.A(net789),
    .B(_01178_),
    .Y(_01305_));
 sky130_fd_sc_hd__a21oi_1 _06179_ (.A1(_01304_),
    .A2(_01305_),
    .B1(net103),
    .Y(_00029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_569 ();
 sky130_fd_sc_hd__nand2_1 _06182_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01171_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_1 _06183_ (.A(net539),
    .B(_01178_),
    .Y(_01309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_568 ();
 sky130_fd_sc_hd__a21oi_1 _06185_ (.A1(_01308_),
    .A2(_01309_),
    .B1(net103),
    .Y(_00030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_566 ();
 sky130_fd_sc_hd__nand2_1 _06188_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_01171_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _06189_ (.A(net1381),
    .B(_01178_),
    .Y(_01314_));
 sky130_fd_sc_hd__a21oi_1 _06190_ (.A1(_01313_),
    .A2(_01314_),
    .B1(net103),
    .Y(_00031_));
 sky130_fd_sc_hd__nand2b_4 _06191_ (.A_N(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .Y(_01315_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_565 ();
 sky130_fd_sc_hd__nand2b_4 _06193_ (.A_N(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .Y(_01317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_564 ();
 sky130_fd_sc_hd__nor3_4 _06195_ (.A(_01162_),
    .B(_01315_),
    .C(_01317_),
    .Y(_01319_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_563 ();
 sky130_fd_sc_hd__nand2_1 _06197_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net89),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_8 _06198_ (.A(_01315_),
    .B(_01317_),
    .Y(_01322_));
 sky130_fd_sc_hd__nand2_8 _06199_ (.A(_01174_),
    .B(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_562 ();
 sky130_fd_sc_hd__nand2_1 _06201_ (.A(net785),
    .B(_01323_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21oi_1 _06202_ (.A1(_01321_),
    .A2(_01325_),
    .B1(net104),
    .Y(_00032_));
 sky130_fd_sc_hd__nand2_1 _06203_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net88),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _06204_ (.A(net456),
    .B(_01323_),
    .Y(_01327_));
 sky130_fd_sc_hd__a21oi_1 _06205_ (.A1(_01326_),
    .A2(_01327_),
    .B1(net107),
    .Y(_00033_));
 sky130_fd_sc_hd__nand2_1 _06206_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net88),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _06207_ (.A(net533),
    .B(_01323_),
    .Y(_01329_));
 sky130_fd_sc_hd__a21oi_1 _06208_ (.A1(_01328_),
    .A2(_01329_),
    .B1(CPU_reset_a4),
    .Y(_00034_));
 sky130_fd_sc_hd__nand2_1 _06209_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net87),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _06210_ (.A(net241),
    .B(_01323_),
    .Y(_01331_));
 sky130_fd_sc_hd__a21oi_1 _06211_ (.A1(_01330_),
    .A2(_01331_),
    .B1(net102),
    .Y(_00035_));
 sky130_fd_sc_hd__nand2_1 _06212_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net87),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _06213_ (.A(net909),
    .B(_01323_),
    .Y(_01333_));
 sky130_fd_sc_hd__a21oi_1 _06214_ (.A1(_01332_),
    .A2(_01333_),
    .B1(net106),
    .Y(_00036_));
 sky130_fd_sc_hd__nand2_1 _06215_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net87),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_1 _06216_ (.A(net229),
    .B(_01323_),
    .Y(_01335_));
 sky130_fd_sc_hd__a21oi_1 _06217_ (.A1(_01334_),
    .A2(_01335_),
    .B1(net107),
    .Y(_00037_));
 sky130_fd_sc_hd__nand2_1 _06218_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net87),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _06219_ (.A(net952),
    .B(_01323_),
    .Y(_01337_));
 sky130_fd_sc_hd__a21oi_1 _06220_ (.A1(_01336_),
    .A2(_01337_),
    .B1(net105),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _06221_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net89),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _06222_ (.A(net942),
    .B(_01323_),
    .Y(_01339_));
 sky130_fd_sc_hd__a21oi_1 _06223_ (.A1(_01338_),
    .A2(_01339_),
    .B1(net105),
    .Y(_00039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_561 ();
 sky130_fd_sc_hd__nand2_1 _06225_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net87),
    .Y(_01341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_560 ();
 sky130_fd_sc_hd__nand2_1 _06227_ (.A(net446),
    .B(_01323_),
    .Y(_01343_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_559 ();
 sky130_fd_sc_hd__a21oi_1 _06229_ (.A1(_01341_),
    .A2(_01343_),
    .B1(net102),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _06230_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net87),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_1 _06231_ (.A(net343),
    .B(_01323_),
    .Y(_01346_));
 sky130_fd_sc_hd__a21oi_1 _06232_ (.A1(_01345_),
    .A2(_01346_),
    .B1(net106),
    .Y(_00041_));
 sky130_fd_sc_hd__nand2_1 _06233_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net87),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _06234_ (.A(net1206),
    .B(_01323_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21oi_1 _06235_ (.A1(_01347_),
    .A2(_01348_),
    .B1(CPU_reset_a4),
    .Y(_00042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_558 ();
 sky130_fd_sc_hd__nand2_1 _06237_ (.A(net1073),
    .B(_01323_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _06238_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01319_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand3b_1 _06239_ (.A_N(net103),
    .B(_01350_),
    .C(_01351_),
    .Y(_00043_));
 sky130_fd_sc_hd__nand2_1 _06240_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net89),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _06241_ (.A(net478),
    .B(_01323_),
    .Y(_01353_));
 sky130_fd_sc_hd__a21oi_1 _06242_ (.A1(_01352_),
    .A2(_01353_),
    .B1(net102),
    .Y(_00044_));
 sky130_fd_sc_hd__nand2_1 _06243_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net87),
    .Y(_01354_));
 sky130_fd_sc_hd__nand2_1 _06244_ (.A(net349),
    .B(_01323_),
    .Y(_01355_));
 sky130_fd_sc_hd__a21oi_1 _06245_ (.A1(_01354_),
    .A2(_01355_),
    .B1(net104),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _06246_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net88),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _06247_ (.A(net1101),
    .B(_01323_),
    .Y(_01357_));
 sky130_fd_sc_hd__a21oi_1 _06248_ (.A1(_01356_),
    .A2(_01357_),
    .B1(CPU_reset_a4),
    .Y(_00046_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net89),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_1 _06250_ (.A(net819),
    .B(_01323_),
    .Y(_01359_));
 sky130_fd_sc_hd__a21oi_1 _06251_ (.A1(_01358_),
    .A2(_01359_),
    .B1(net102),
    .Y(_00047_));
 sky130_fd_sc_hd__nand2_1 _06252_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net87),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _06253_ (.A(net555),
    .B(_01323_),
    .Y(_01361_));
 sky130_fd_sc_hd__a21oi_1 _06254_ (.A1(_01360_),
    .A2(_01361_),
    .B1(CPU_reset_a4),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _06255_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net87),
    .Y(_01362_));
 sky130_fd_sc_hd__nand2_1 _06256_ (.A(net480),
    .B(_01323_),
    .Y(_01363_));
 sky130_fd_sc_hd__a21oi_1 _06257_ (.A1(_01362_),
    .A2(_01363_),
    .B1(net106),
    .Y(_00049_));
 sky130_fd_sc_hd__nand2_1 _06258_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net88),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _06259_ (.A(net946),
    .B(_01323_),
    .Y(_01365_));
 sky130_fd_sc_hd__a21oi_1 _06260_ (.A1(_01364_),
    .A2(_01365_),
    .B1(CPU_reset_a4),
    .Y(_00050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_557 ();
 sky130_fd_sc_hd__nand2_1 _06262_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net88),
    .Y(_01367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_556 ();
 sky130_fd_sc_hd__nand2_1 _06264_ (.A(net850),
    .B(_01323_),
    .Y(_01369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_555 ();
 sky130_fd_sc_hd__a21oi_1 _06266_ (.A1(_01367_),
    .A2(_01369_),
    .B1(net105),
    .Y(_00051_));
 sky130_fd_sc_hd__nand2_1 _06267_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net87),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2_1 _06268_ (.A(net984),
    .B(_01323_),
    .Y(_01372_));
 sky130_fd_sc_hd__a21oi_1 _06269_ (.A1(_01371_),
    .A2(_01372_),
    .B1(net102),
    .Y(_00052_));
 sky130_fd_sc_hd__nand2_1 _06270_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net87),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _06271_ (.A(net585),
    .B(_01323_),
    .Y(_01374_));
 sky130_fd_sc_hd__a21oi_1 _06272_ (.A1(_01373_),
    .A2(_01374_),
    .B1(net107),
    .Y(_00053_));
 sky130_fd_sc_hd__nand2_1 _06273_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01319_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _06274_ (.A(net466),
    .B(_01323_),
    .Y(_01376_));
 sky130_fd_sc_hd__a21oi_1 _06275_ (.A1(_01375_),
    .A2(_01376_),
    .B1(net103),
    .Y(_00054_));
 sky130_fd_sc_hd__nand2_1 _06276_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net88),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _06277_ (.A(net482),
    .B(_01323_),
    .Y(_01378_));
 sky130_fd_sc_hd__a21oi_1 _06278_ (.A1(_01377_),
    .A2(_01378_),
    .B1(net107),
    .Y(_00055_));
 sky130_fd_sc_hd__nand2_1 _06279_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net88),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _06280_ (.A(net903),
    .B(_01323_),
    .Y(_01380_));
 sky130_fd_sc_hd__a21oi_1 _06281_ (.A1(_01379_),
    .A2(_01380_),
    .B1(net105),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _06282_ (.A(net1127),
    .B(_01323_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _06283_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01319_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand3b_1 _06284_ (.A_N(net103),
    .B(_01381_),
    .C(_01382_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_1 _06285_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net89),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2_1 _06286_ (.A(net920),
    .B(_01323_),
    .Y(_01384_));
 sky130_fd_sc_hd__a21oi_1 _06287_ (.A1(_01383_),
    .A2(_01384_),
    .B1(net104),
    .Y(_00058_));
 sky130_fd_sc_hd__nand2_1 _06288_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01319_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(net361),
    .B(_01323_),
    .Y(_01386_));
 sky130_fd_sc_hd__a21oi_1 _06290_ (.A1(_01385_),
    .A2(_01386_),
    .B1(net105),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _06291_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net88),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _06292_ (.A(net950),
    .B(_01323_),
    .Y(_01388_));
 sky130_fd_sc_hd__a21oi_1 _06293_ (.A1(_01387_),
    .A2(_01388_),
    .B1(net107),
    .Y(_00060_));
 sky130_fd_sc_hd__nand2_1 _06294_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net89),
    .Y(_01389_));
 sky130_fd_sc_hd__nand2_1 _06295_ (.A(net1034),
    .B(_01323_),
    .Y(_01390_));
 sky130_fd_sc_hd__a21oi_1 _06296_ (.A1(_01389_),
    .A2(_01390_),
    .B1(net104),
    .Y(_00061_));
 sky130_fd_sc_hd__nand2_1 _06297_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01319_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _06298_ (.A(net492),
    .B(_01323_),
    .Y(_01392_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_554 ();
 sky130_fd_sc_hd__a21oi_1 _06300_ (.A1(_01391_),
    .A2(_01392_),
    .B1(net103),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _06301_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net89),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _06302_ (.A(net454),
    .B(_01323_),
    .Y(_01395_));
 sky130_fd_sc_hd__a21oi_1 _06303_ (.A1(_01394_),
    .A2(_01395_),
    .B1(net105),
    .Y(_00063_));
 sky130_fd_sc_hd__nand2_8 _06304_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_8 _06305_ (.A(_01317_),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_8 _06306_ (.A(_01174_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_553 ();
 sky130_fd_sc_hd__nand2_1 _06308_ (.A(net980),
    .B(_01398_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor3_4 _06309_ (.A(_01162_),
    .B(_01317_),
    .C(_01396_),
    .Y(_01401_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_552 ();
 sky130_fd_sc_hd__nand2_1 _06311_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(_01401_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3b_1 _06312_ (.A_N(net104),
    .B(_01400_),
    .C(_01403_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand2_1 _06313_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net86),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(net393),
    .B(_01398_),
    .Y(_01405_));
 sky130_fd_sc_hd__a21oi_1 _06315_ (.A1(_01404_),
    .A2(_01405_),
    .B1(net105),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_1 _06316_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net86),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _06317_ (.A(net614),
    .B(_01398_),
    .Y(_01407_));
 sky130_fd_sc_hd__a21oi_1 _06318_ (.A1(_01406_),
    .A2(_01407_),
    .B1(CPU_reset_a4),
    .Y(_00066_));
 sky130_fd_sc_hd__nand2_1 _06319_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(_01401_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _06320_ (.A(net355),
    .B(_01398_),
    .Y(_01409_));
 sky130_fd_sc_hd__a21oi_1 _06321_ (.A1(_01408_),
    .A2(_01409_),
    .B1(net102),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net85),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_1 _06323_ (.A(net347),
    .B(_01398_),
    .Y(_01411_));
 sky130_fd_sc_hd__a21oi_1 _06324_ (.A1(_01410_),
    .A2(_01411_),
    .B1(net106),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net85),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(net866),
    .B(_01398_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21oi_1 _06327_ (.A1(_01412_),
    .A2(_01413_),
    .B1(net107),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_1 _06328_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net85),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _06329_ (.A(net632),
    .B(_01398_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21oi_1 _06330_ (.A1(_01414_),
    .A2(_01415_),
    .B1(net102),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _06331_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net86),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2_1 _06332_ (.A(net978),
    .B(_01398_),
    .Y(_01417_));
 sky130_fd_sc_hd__a21oi_1 _06333_ (.A1(_01416_),
    .A2(_01417_),
    .B1(net105),
    .Y(_00071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_551 ();
 sky130_fd_sc_hd__nand2_1 _06335_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(_01401_),
    .Y(_01419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_550 ();
 sky130_fd_sc_hd__nand2_1 _06337_ (.A(net529),
    .B(_01398_),
    .Y(_01421_));
 sky130_fd_sc_hd__a21oi_1 _06338_ (.A1(_01419_),
    .A2(_01421_),
    .B1(net102),
    .Y(_00072_));
 sky130_fd_sc_hd__nand2_1 _06339_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net85),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _06340_ (.A(net602),
    .B(_01398_),
    .Y(_01423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_549 ();
 sky130_fd_sc_hd__a21oi_1 _06342_ (.A1(_01422_),
    .A2(_01423_),
    .B1(net106),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_1 _06343_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net85),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _06344_ (.A(net411),
    .B(_01398_),
    .Y(_01426_));
 sky130_fd_sc_hd__a21oi_1 _06345_ (.A1(_01425_),
    .A2(_01426_),
    .B1(net106),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_1 _06346_ (.A(net1208),
    .B(_01398_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _06347_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01401_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand3b_1 _06348_ (.A_N(net103),
    .B(_01427_),
    .C(_01428_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand2_1 _06349_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(_01401_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _06350_ (.A(net335),
    .B(_01398_),
    .Y(_01430_));
 sky130_fd_sc_hd__a21oi_1 _06351_ (.A1(_01429_),
    .A2(_01430_),
    .B1(net102),
    .Y(_00076_));
 sky130_fd_sc_hd__nand2_1 _06352_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net85),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _06353_ (.A(net680),
    .B(_01398_),
    .Y(_01432_));
 sky130_fd_sc_hd__a21oi_1 _06354_ (.A1(_01431_),
    .A2(_01432_),
    .B1(net104),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net86),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _06356_ (.A(net1022),
    .B(_01398_),
    .Y(_01434_));
 sky130_fd_sc_hd__a21oi_1 _06357_ (.A1(_01433_),
    .A2(_01434_),
    .B1(CPU_reset_a4),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_1 _06358_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_01401_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(net884),
    .B(_01398_),
    .Y(_01436_));
 sky130_fd_sc_hd__a21oi_1 _06360_ (.A1(_01435_),
    .A2(_01436_),
    .B1(net104),
    .Y(_00079_));
 sky130_fd_sc_hd__nand2_1 _06361_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net86),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _06362_ (.A(net1008),
    .B(_01398_),
    .Y(_01438_));
 sky130_fd_sc_hd__a21oi_1 _06363_ (.A1(_01437_),
    .A2(_01438_),
    .B1(CPU_reset_a4),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_1 _06364_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net85),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _06365_ (.A(net1057),
    .B(_01398_),
    .Y(_01440_));
 sky130_fd_sc_hd__a21oi_1 _06366_ (.A1(_01439_),
    .A2(_01440_),
    .B1(net106),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _06367_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net86),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _06368_ (.A(net940),
    .B(_01398_),
    .Y(_01442_));
 sky130_fd_sc_hd__a21oi_1 _06369_ (.A1(_01441_),
    .A2(_01442_),
    .B1(net106),
    .Y(_00082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_548 ();
 sky130_fd_sc_hd__nand2_1 _06371_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net85),
    .Y(_01444_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_547 ();
 sky130_fd_sc_hd__nand2_1 _06373_ (.A(net896),
    .B(_01398_),
    .Y(_01446_));
 sky130_fd_sc_hd__a21oi_1 _06374_ (.A1(_01444_),
    .A2(_01446_),
    .B1(net105),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _06375_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net85),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _06376_ (.A(net442),
    .B(_01398_),
    .Y(_01448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_545 ();
 sky130_fd_sc_hd__a21oi_1 _06379_ (.A1(_01447_),
    .A2(_01448_),
    .B1(net104),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net85),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _06381_ (.A(net559),
    .B(_01398_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21oi_1 _06382_ (.A1(_01451_),
    .A2(_01452_),
    .B1(net107),
    .Y(_00085_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01401_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _06384_ (.A(net805),
    .B(_01398_),
    .Y(_01454_));
 sky130_fd_sc_hd__a21oi_1 _06385_ (.A1(_01453_),
    .A2(_01454_),
    .B1(net103),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _06386_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net86),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _06387_ (.A(net407),
    .B(_01398_),
    .Y(_01456_));
 sky130_fd_sc_hd__a21oi_1 _06388_ (.A1(_01455_),
    .A2(_01456_),
    .B1(net107),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_1 _06389_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net86),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(net620),
    .B(_01398_),
    .Y(_01458_));
 sky130_fd_sc_hd__a21oi_1 _06391_ (.A1(_01457_),
    .A2(_01458_),
    .B1(net105),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_1 _06392_ (.A(net1059),
    .B(_01398_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_1 _06393_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01401_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand3b_1 _06394_ (.A_N(net103),
    .B(_01459_),
    .C(_01460_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_01401_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _06396_ (.A(net745),
    .B(_01398_),
    .Y(_01462_));
 sky130_fd_sc_hd__a21oi_1 _06397_ (.A1(_01461_),
    .A2(_01462_),
    .B1(net104),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_1 _06398_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(net86),
    .Y(_01463_));
 sky130_fd_sc_hd__nand2_1 _06399_ (.A(net1174),
    .B(_01398_),
    .Y(_01464_));
 sky130_fd_sc_hd__a21oi_1 _06400_ (.A1(_01463_),
    .A2(_01464_),
    .B1(net105),
    .Y(_00091_));
 sky130_fd_sc_hd__nand2_1 _06401_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net86),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _06402_ (.A(net630),
    .B(_01398_),
    .Y(_01466_));
 sky130_fd_sc_hd__a21oi_1 _06403_ (.A1(_01465_),
    .A2(_01466_),
    .B1(CPU_reset_a4),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_1 _06404_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_01401_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _06405_ (.A(net968),
    .B(_01398_),
    .Y(_01468_));
 sky130_fd_sc_hd__a21oi_1 _06406_ (.A1(_01467_),
    .A2(_01468_),
    .B1(net103),
    .Y(_00093_));
 sky130_fd_sc_hd__nand2_1 _06407_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01401_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _06408_ (.A(net672),
    .B(_01398_),
    .Y(_01470_));
 sky130_fd_sc_hd__a21oi_1 _06409_ (.A1(_01469_),
    .A2(_01470_),
    .B1(net103),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_1 _06410_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_01401_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _06411_ (.A(net1329),
    .B(_01398_),
    .Y(_01472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_544 ();
 sky130_fd_sc_hd__a21oi_1 _06413_ (.A1(_01471_),
    .A2(_01472_),
    .B1(net103),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_8 _06414_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .Y(_01474_));
 sky130_fd_sc_hd__nor4_4 _06415_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_01162_),
    .D(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_543 ();
 sky130_fd_sc_hd__nand2_1 _06417_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net84),
    .Y(_01477_));
 sky130_fd_sc_hd__nor3_4 _06418_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_01474_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_8 _06419_ (.A(_01174_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_542 ();
 sky130_fd_sc_hd__nand2_1 _06421_ (.A(net551),
    .B(_01479_),
    .Y(_01481_));
 sky130_fd_sc_hd__a21oi_1 _06422_ (.A1(_01477_),
    .A2(_01481_),
    .B1(net104),
    .Y(_00096_));
 sky130_fd_sc_hd__nand2_1 _06423_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net83),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _06424_ (.A(net437),
    .B(_01479_),
    .Y(_01483_));
 sky130_fd_sc_hd__a21oi_1 _06425_ (.A1(_01482_),
    .A2(_01483_),
    .B1(net105),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net82),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(net834),
    .B(_01479_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21oi_1 _06428_ (.A1(_01484_),
    .A2(_01485_),
    .B1(CPU_reset_a4),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _06429_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net84),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _06430_ (.A(net1105),
    .B(_01479_),
    .Y(_01487_));
 sky130_fd_sc_hd__a21oi_1 _06431_ (.A1(_01486_),
    .A2(_01487_),
    .B1(net107),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2_1 _06432_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net83),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(net329),
    .B(_01479_),
    .Y(_01489_));
 sky130_fd_sc_hd__a21oi_1 _06434_ (.A1(_01488_),
    .A2(_01489_),
    .B1(net106),
    .Y(_00100_));
 sky130_fd_sc_hd__nand2_1 _06435_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net83),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _06436_ (.A(net557),
    .B(_01479_),
    .Y(_01491_));
 sky130_fd_sc_hd__a21oi_1 _06437_ (.A1(_01490_),
    .A2(_01491_),
    .B1(net106),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net84),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _06439_ (.A(net1121),
    .B(_01479_),
    .Y(_01493_));
 sky130_fd_sc_hd__a21oi_1 _06440_ (.A1(_01492_),
    .A2(_01493_),
    .B1(net102),
    .Y(_00102_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net84),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _06442_ (.A(net801),
    .B(_01479_),
    .Y(_01495_));
 sky130_fd_sc_hd__a21oi_1 _06443_ (.A1(_01494_),
    .A2(_01495_),
    .B1(net104),
    .Y(_00103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_541 ();
 sky130_fd_sc_hd__nand2_1 _06445_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net84),
    .Y(_01497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_540 ();
 sky130_fd_sc_hd__nand2_1 _06447_ (.A(net460),
    .B(_01479_),
    .Y(_01499_));
 sky130_fd_sc_hd__a21oi_1 _06448_ (.A1(_01497_),
    .A2(_01499_),
    .B1(net102),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _06449_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net83),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _06450_ (.A(net700),
    .B(_01479_),
    .Y(_01501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_539 ();
 sky130_fd_sc_hd__a21oi_1 _06452_ (.A1(_01500_),
    .A2(_01501_),
    .B1(net106),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_1 _06453_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net82),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _06454_ (.A(net409),
    .B(_01479_),
    .Y(_01504_));
 sky130_fd_sc_hd__a21oi_1 _06455_ (.A1(_01503_),
    .A2(_01504_),
    .B1(CPU_reset_a4),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _06456_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01475_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _06457_ (.A(net787),
    .B(_01479_),
    .Y(_01506_));
 sky130_fd_sc_hd__a21oi_1 _06458_ (.A1(_01505_),
    .A2(_01506_),
    .B1(net103),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _06459_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net84),
    .Y(_01507_));
 sky130_fd_sc_hd__nand2_1 _06460_ (.A(net624),
    .B(_01479_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21oi_1 _06461_ (.A1(_01507_),
    .A2(_01508_),
    .B1(net102),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net84),
    .Y(_01509_));
 sky130_fd_sc_hd__nand2_1 _06463_ (.A(net476),
    .B(_01479_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21oi_1 _06464_ (.A1(_01509_),
    .A2(_01510_),
    .B1(net104),
    .Y(_00109_));
 sky130_fd_sc_hd__nand2_1 _06465_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net82),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _06466_ (.A(net856),
    .B(_01479_),
    .Y(_01512_));
 sky130_fd_sc_hd__a21oi_1 _06467_ (.A1(_01511_),
    .A2(_01512_),
    .B1(CPU_reset_a4),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _06468_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_01475_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _06469_ (.A(net922),
    .B(_01479_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_1 _06470_ (.A1(_01513_),
    .A2(_01514_),
    .B1(net102),
    .Y(_00111_));
 sky130_fd_sc_hd__nand2_1 _06471_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net82),
    .Y(_01515_));
 sky130_fd_sc_hd__nand2_1 _06472_ (.A(net1109),
    .B(_01479_),
    .Y(_01516_));
 sky130_fd_sc_hd__a21oi_1 _06473_ (.A1(_01515_),
    .A2(_01516_),
    .B1(CPU_reset_a4),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net83),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _06475_ (.A(net253),
    .B(_01479_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21oi_1 _06476_ (.A1(_01517_),
    .A2(_01518_),
    .B1(net106),
    .Y(_00113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_538 ();
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net82),
    .Y(_01520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_537 ();
 sky130_fd_sc_hd__nand2_1 _06480_ (.A(net880),
    .B(_01479_),
    .Y(_01522_));
 sky130_fd_sc_hd__a21oi_1 _06481_ (.A1(_01520_),
    .A2(_01522_),
    .B1(net106),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _06482_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net83),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _06483_ (.A(net452),
    .B(_01479_),
    .Y(_01524_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_536 ();
 sky130_fd_sc_hd__a21oi_1 _06485_ (.A1(_01523_),
    .A2(_01524_),
    .B1(net105),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _06486_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net83),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _06487_ (.A(net823),
    .B(_01479_),
    .Y(_01527_));
 sky130_fd_sc_hd__a21oi_1 _06488_ (.A1(_01526_),
    .A2(_01527_),
    .B1(net107),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_1 _06489_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net83),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _06490_ (.A(net779),
    .B(_01479_),
    .Y(_01529_));
 sky130_fd_sc_hd__a21oi_1 _06491_ (.A1(_01528_),
    .A2(_01529_),
    .B1(net107),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _06492_ (.A(net1219),
    .B(_01479_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01475_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand3b_1 _06494_ (.A_N(net103),
    .B(_01530_),
    .C(_01531_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net82),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _06496_ (.A(net682),
    .B(_01479_),
    .Y(_01533_));
 sky130_fd_sc_hd__a21oi_1 _06497_ (.A1(_01532_),
    .A2(_01533_),
    .B1(net106),
    .Y(_00119_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net84),
    .Y(_01534_));
 sky130_fd_sc_hd__nand2_1 _06499_ (.A(net1533),
    .B(_01479_),
    .Y(_01535_));
 sky130_fd_sc_hd__a21oi_1 _06500_ (.A1(_01534_),
    .A2(_01535_),
    .B1(net105),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _06501_ (.A(net1231),
    .B(_01479_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _06502_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01475_),
    .Y(_01537_));
 sky130_fd_sc_hd__nand3b_1 _06503_ (.A_N(net103),
    .B(_01536_),
    .C(_01537_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_1 _06504_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_01475_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand2_1 _06505_ (.A(net517),
    .B(_01479_),
    .Y(_01539_));
 sky130_fd_sc_hd__a21oi_1 _06506_ (.A1(_01538_),
    .A2(_01539_),
    .B1(net104),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _06507_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01475_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _06508_ (.A(net1344),
    .B(_01479_),
    .Y(_01541_));
 sky130_fd_sc_hd__a21oi_1 _06509_ (.A1(_01540_),
    .A2(_01541_),
    .B1(net105),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _06510_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net82),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _06511_ (.A(net1202),
    .B(_01479_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21oi_1 _06512_ (.A1(_01542_),
    .A2(_01543_),
    .B1(CPU_reset_a4),
    .Y(_00124_));
 sky130_fd_sc_hd__nand2_1 _06513_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_01475_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(net628),
    .B(_01479_),
    .Y(_01545_));
 sky130_fd_sc_hd__a21oi_1 _06515_ (.A1(_01544_),
    .A2(_01545_),
    .B1(net103),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _06516_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01475_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _06517_ (.A(net761),
    .B(_01479_),
    .Y(_01547_));
 sky130_fd_sc_hd__a21oi_1 _06518_ (.A1(_01546_),
    .A2(_01547_),
    .B1(net103),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _06519_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net84),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _06520_ (.A(net1193),
    .B(_01479_),
    .Y(_01549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_535 ();
 sky130_fd_sc_hd__a21oi_1 _06522_ (.A1(_01548_),
    .A2(_01549_),
    .B1(net104),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2b_4 _06523_ (.A_N(\CPU_dmem_addr_a4[1] ),
    .B(\CPU_dmem_addr_a4[0] ),
    .Y(_01551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_534 ();
 sky130_fd_sc_hd__nor2_8 _06525_ (.A(_01474_),
    .B(_01551_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_8 _06526_ (.A(_01174_),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_533 ();
 sky130_fd_sc_hd__nand2_1 _06528_ (.A(net1251),
    .B(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor3_4 _06529_ (.A(_01162_),
    .B(_01474_),
    .C(_01551_),
    .Y(_01557_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_532 ();
 sky130_fd_sc_hd__nand2_1 _06531_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net78),
    .Y(_01559_));
 sky130_fd_sc_hd__nand3b_1 _06532_ (.A_N(net104),
    .B(_01556_),
    .C(_01559_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _06533_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net79),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(net1129),
    .B(_01554_),
    .Y(_01561_));
 sky130_fd_sc_hd__a21oi_1 _06535_ (.A1(_01560_),
    .A2(_01561_),
    .B1(net105),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net79),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _06537_ (.A(net670),
    .B(_01554_),
    .Y(_01563_));
 sky130_fd_sc_hd__a21oi_1 _06538_ (.A1(_01562_),
    .A2(_01563_),
    .B1(CPU_reset_a4),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _06539_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net78),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _06540_ (.A(net458),
    .B(_01554_),
    .Y(_01565_));
 sky130_fd_sc_hd__a21oi_1 _06541_ (.A1(_01564_),
    .A2(_01565_),
    .B1(net107),
    .Y(_00131_));
 sky130_fd_sc_hd__nand2_1 _06542_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net79),
    .Y(_01566_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(net1111),
    .B(_01554_),
    .Y(_01567_));
 sky130_fd_sc_hd__a21oi_1 _06544_ (.A1(_01566_),
    .A2(_01567_),
    .B1(net106),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _06545_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net79),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(net249),
    .B(_01554_),
    .Y(_01569_));
 sky130_fd_sc_hd__a21oi_1 _06547_ (.A1(_01568_),
    .A2(_01569_),
    .B1(net107),
    .Y(_00133_));
 sky130_fd_sc_hd__nand2_1 _06548_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net79),
    .Y(_01570_));
 sky130_fd_sc_hd__nand2_1 _06549_ (.A(net694),
    .B(_01554_),
    .Y(_01571_));
 sky130_fd_sc_hd__a21oi_1 _06550_ (.A1(_01570_),
    .A2(_01571_),
    .B1(net104),
    .Y(_00134_));
 sky130_fd_sc_hd__nand2_1 _06551_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(_01557_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _06552_ (.A(net711),
    .B(_01554_),
    .Y(_01573_));
 sky130_fd_sc_hd__a21oi_1 _06553_ (.A1(_01572_),
    .A2(_01573_),
    .B1(net105),
    .Y(_00135_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_531 ();
 sky130_fd_sc_hd__nand2_1 _06555_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net78),
    .Y(_01575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_530 ();
 sky130_fd_sc_hd__nand2_1 _06557_ (.A(net656),
    .B(_01554_),
    .Y(_01577_));
 sky130_fd_sc_hd__a21oi_1 _06558_ (.A1(_01575_),
    .A2(_01577_),
    .B1(net102),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_1 _06559_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net79),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _06560_ (.A(net737),
    .B(_01554_),
    .Y(_01579_));
 sky130_fd_sc_hd__a21oi_1 _06561_ (.A1(_01578_),
    .A2(_01579_),
    .B1(net106),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _06562_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net79),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_1 _06563_ (.A(net341),
    .B(_01554_),
    .Y(_01581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_529 ();
 sky130_fd_sc_hd__a21oi_1 _06565_ (.A1(_01580_),
    .A2(_01581_),
    .B1(CPU_reset_a4),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01557_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _06567_ (.A(net505),
    .B(_01554_),
    .Y(_01584_));
 sky130_fd_sc_hd__a21oi_1 _06568_ (.A1(_01583_),
    .A2(_01584_),
    .B1(net103),
    .Y(_00139_));
 sky130_fd_sc_hd__nand2_1 _06569_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net78),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _06570_ (.A(net1147),
    .B(_01554_),
    .Y(_01586_));
 sky130_fd_sc_hd__a21oi_1 _06571_ (.A1(_01585_),
    .A2(_01586_),
    .B1(net102),
    .Y(_00140_));
 sky130_fd_sc_hd__nand2_1 _06572_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net78),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _06573_ (.A(net876),
    .B(_01554_),
    .Y(_01588_));
 sky130_fd_sc_hd__a21oi_1 _06574_ (.A1(_01587_),
    .A2(_01588_),
    .B1(net104),
    .Y(_00141_));
 sky130_fd_sc_hd__nand2_1 _06575_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net79),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_1 _06576_ (.A(net809),
    .B(_01554_),
    .Y(_01590_));
 sky130_fd_sc_hd__a21oi_1 _06577_ (.A1(_01589_),
    .A2(_01590_),
    .B1(CPU_reset_a4),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net78),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _06579_ (.A(net901),
    .B(_01554_),
    .Y(_01592_));
 sky130_fd_sc_hd__a21oi_1 _06580_ (.A1(_01591_),
    .A2(_01592_),
    .B1(net104),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _06581_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net79),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _06582_ (.A(net1093),
    .B(_01554_),
    .Y(_01594_));
 sky130_fd_sc_hd__a21oi_1 _06583_ (.A1(_01593_),
    .A2(_01594_),
    .B1(CPU_reset_a4),
    .Y(_00144_));
 sky130_fd_sc_hd__nand2_1 _06584_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net79),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_1 _06585_ (.A(net365),
    .B(_01554_),
    .Y(_01596_));
 sky130_fd_sc_hd__a21oi_1 _06586_ (.A1(_01595_),
    .A2(_01596_),
    .B1(net106),
    .Y(_00145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_528 ();
 sky130_fd_sc_hd__nand2_1 _06588_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net79),
    .Y(_01598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_527 ();
 sky130_fd_sc_hd__nand2_1 _06590_ (.A(net431),
    .B(_01554_),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_1 _06591_ (.A1(_01598_),
    .A2(_01600_),
    .B1(CPU_reset_a4),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_1 _06592_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net79),
    .Y(_01601_));
 sky130_fd_sc_hd__nand2_1 _06593_ (.A(net815),
    .B(_01554_),
    .Y(_01602_));
 sky130_fd_sc_hd__a21oi_1 _06594_ (.A1(_01601_),
    .A2(_01602_),
    .B1(net105),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _06595_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net79),
    .Y(_01603_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(net1014),
    .B(_01554_),
    .Y(_01604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_526 ();
 sky130_fd_sc_hd__a21oi_1 _06598_ (.A1(_01603_),
    .A2(_01604_),
    .B1(net104),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _06599_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net78),
    .Y(_01606_));
 sky130_fd_sc_hd__nand2_1 _06600_ (.A(net813),
    .B(_01554_),
    .Y(_01607_));
 sky130_fd_sc_hd__a21oi_1 _06601_ (.A1(_01606_),
    .A2(_01607_),
    .B1(net107),
    .Y(_00149_));
 sky130_fd_sc_hd__nand2_1 _06602_ (.A(net1348),
    .B(_01554_),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2_1 _06603_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01557_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand3b_1 _06604_ (.A_N(net103),
    .B(_01608_),
    .C(_01609_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2_1 _06605_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net79),
    .Y(_01610_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(net1046),
    .B(_01554_),
    .Y(_01611_));
 sky130_fd_sc_hd__a21oi_1 _06607_ (.A1(_01610_),
    .A2(_01611_),
    .B1(net106),
    .Y(_00151_));
 sky130_fd_sc_hd__nand2_1 _06608_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(_01557_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand2_1 _06609_ (.A(net913),
    .B(_01554_),
    .Y(_01613_));
 sky130_fd_sc_hd__a21oi_1 _06610_ (.A1(_01612_),
    .A2(_01613_),
    .B1(net105),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _06611_ (.A(net1264),
    .B(_01554_),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_1 _06612_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01557_),
    .Y(_01615_));
 sky130_fd_sc_hd__nand3b_1 _06613_ (.A_N(net103),
    .B(_01614_),
    .C(_01615_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _06614_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net78),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _06615_ (.A(net654),
    .B(_01554_),
    .Y(_01617_));
 sky130_fd_sc_hd__a21oi_1 _06616_ (.A1(_01616_),
    .A2(_01617_),
    .B1(net103),
    .Y(_00154_));
 sky130_fd_sc_hd__nand2_1 _06617_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01557_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(net994),
    .B(_01554_),
    .Y(_01619_));
 sky130_fd_sc_hd__a21oi_1 _06619_ (.A1(_01618_),
    .A2(_01619_),
    .B1(net105),
    .Y(_00155_));
 sky130_fd_sc_hd__nand2_1 _06620_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net79),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _06621_ (.A(net291),
    .B(_01554_),
    .Y(_01621_));
 sky130_fd_sc_hd__a21oi_1 _06622_ (.A1(_01620_),
    .A2(_01621_),
    .B1(CPU_reset_a4),
    .Y(_00156_));
 sky130_fd_sc_hd__nand2_1 _06623_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net78),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _06624_ (.A(net678),
    .B(_01554_),
    .Y(_01623_));
 sky130_fd_sc_hd__a21oi_1 _06625_ (.A1(_01622_),
    .A2(_01623_),
    .B1(net103),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _06626_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01557_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _06627_ (.A(net1152),
    .B(_01554_),
    .Y(_01625_));
 sky130_fd_sc_hd__a21oi_1 _06628_ (.A1(_01624_),
    .A2(_01625_),
    .B1(net103),
    .Y(_00158_));
 sky130_fd_sc_hd__nand2_1 _06629_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net78),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _06630_ (.A(net1246),
    .B(_01554_),
    .Y(_01627_));
 sky130_fd_sc_hd__a21oi_1 _06631_ (.A1(_01626_),
    .A2(_01627_),
    .B1(net103),
    .Y(_00159_));
 sky130_fd_sc_hd__nor3_4 _06632_ (.A(_01162_),
    .B(_01315_),
    .C(_01474_),
    .Y(_01628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_525 ();
 sky130_fd_sc_hd__nand2_1 _06634_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net77),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_8 _06635_ (.A(_01315_),
    .B(_01474_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand2_8 _06636_ (.A(_01174_),
    .B(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_524 ();
 sky130_fd_sc_hd__nand2_1 _06638_ (.A(net519),
    .B(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_523 ();
 sky130_fd_sc_hd__a21oi_1 _06640_ (.A1(_01630_),
    .A2(_01634_),
    .B1(net104),
    .Y(_00160_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net77),
    .Y(_01636_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(net351),
    .B(_01632_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21oi_1 _06643_ (.A1(_01636_),
    .A2(_01637_),
    .B1(net105),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net76),
    .Y(_01638_));
 sky130_fd_sc_hd__nand2_1 _06645_ (.A(net783),
    .B(_01632_),
    .Y(_01639_));
 sky130_fd_sc_hd__a21oi_1 _06646_ (.A1(_01638_),
    .A2(_01639_),
    .B1(net106),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _06647_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net76),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_1 _06648_ (.A(net777),
    .B(_01632_),
    .Y(_01641_));
 sky130_fd_sc_hd__a21oi_1 _06649_ (.A1(_01640_),
    .A2(_01641_),
    .B1(net102),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net76),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_1 _06651_ (.A(net606),
    .B(_01632_),
    .Y(_01643_));
 sky130_fd_sc_hd__a21oi_1 _06652_ (.A1(_01642_),
    .A2(_01643_),
    .B1(net106),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _06653_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net76),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _06654_ (.A(net964),
    .B(_01632_),
    .Y(_01645_));
 sky130_fd_sc_hd__a21oi_1 _06655_ (.A1(_01644_),
    .A2(_01645_),
    .B1(net107),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _06656_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net77),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _06657_ (.A(net515),
    .B(_01632_),
    .Y(_01647_));
 sky130_fd_sc_hd__a21oi_1 _06658_ (.A1(_01646_),
    .A2(_01647_),
    .B1(net105),
    .Y(_00166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_522 ();
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net77),
    .Y(_01649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_521 ();
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(net1087),
    .B(_01632_),
    .Y(_01651_));
 sky130_fd_sc_hd__a21oi_1 _06663_ (.A1(_01649_),
    .A2(_01651_),
    .B1(net104),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _06664_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net76),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(net275),
    .B(_01632_),
    .Y(_01653_));
 sky130_fd_sc_hd__a21oi_1 _06666_ (.A1(_01652_),
    .A2(_01653_),
    .B1(net102),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _06667_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net76),
    .Y(_01654_));
 sky130_fd_sc_hd__nand2_1 _06668_ (.A(net696),
    .B(_01632_),
    .Y(_01655_));
 sky130_fd_sc_hd__a21oi_1 _06669_ (.A1(_01654_),
    .A2(_01655_),
    .B1(net106),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_1 _06670_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net76),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _06671_ (.A(net357),
    .B(_01632_),
    .Y(_01657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_520 ();
 sky130_fd_sc_hd__a21oi_1 _06673_ (.A1(_01656_),
    .A2(_01657_),
    .B1(CPU_reset_a4),
    .Y(_00170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_519 ();
 sky130_fd_sc_hd__nand2_1 _06675_ (.A(net1300),
    .B(_01632_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _06676_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01628_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand3b_1 _06677_ (.A_N(net103),
    .B(_01660_),
    .C(_01661_),
    .Y(_00171_));
 sky130_fd_sc_hd__nand2_1 _06678_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(_01628_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _06679_ (.A(net1061),
    .B(_01632_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21oi_1 _06680_ (.A1(_01662_),
    .A2(_01663_),
    .B1(net102),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net76),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _06682_ (.A(net575),
    .B(_01632_),
    .Y(_01665_));
 sky130_fd_sc_hd__a21oi_1 _06683_ (.A1(_01664_),
    .A2(_01665_),
    .B1(net104),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _06684_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net76),
    .Y(_01666_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(net227),
    .B(_01632_),
    .Y(_01667_));
 sky130_fd_sc_hd__a21oi_1 _06686_ (.A1(_01666_),
    .A2(_01667_),
    .B1(CPU_reset_a4),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _06687_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_01628_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _06688_ (.A(net664),
    .B(_01632_),
    .Y(_01669_));
 sky130_fd_sc_hd__a21oi_1 _06689_ (.A1(_01668_),
    .A2(_01669_),
    .B1(net102),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _06690_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net76),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(net781),
    .B(_01632_),
    .Y(_01671_));
 sky130_fd_sc_hd__a21oi_1 _06692_ (.A1(_01670_),
    .A2(_01671_),
    .B1(CPU_reset_a4),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _06693_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net76),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_1 _06694_ (.A(net1012),
    .B(_01632_),
    .Y(_01673_));
 sky130_fd_sc_hd__a21oi_1 _06695_ (.A1(_01672_),
    .A2(_01673_),
    .B1(net106),
    .Y(_00177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_518 ();
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net76),
    .Y(_01675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_517 ();
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(net257),
    .B(_01632_),
    .Y(_01677_));
 sky130_fd_sc_hd__a21oi_1 _06700_ (.A1(_01675_),
    .A2(_01677_),
    .B1(net106),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _06701_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net77),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _06702_ (.A(net589),
    .B(_01632_),
    .Y(_01679_));
 sky130_fd_sc_hd__a21oi_1 _06703_ (.A1(_01678_),
    .A2(_01679_),
    .B1(net105),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net76),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _06705_ (.A(net713),
    .B(_01632_),
    .Y(_01681_));
 sky130_fd_sc_hd__a21oi_1 _06706_ (.A1(_01680_),
    .A2(_01681_),
    .B1(net104),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net76),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _06708_ (.A(net541),
    .B(_01632_),
    .Y(_01683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_516 ();
 sky130_fd_sc_hd__a21oi_1 _06710_ (.A1(_01682_),
    .A2(_01683_),
    .B1(net107),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _06711_ (.A(net1221),
    .B(_01632_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _06712_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01628_),
    .Y(_01686_));
 sky130_fd_sc_hd__nand3b_1 _06713_ (.A_N(net103),
    .B(_01685_),
    .C(_01686_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net77),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(net996),
    .B(_01632_),
    .Y(_01688_));
 sky130_fd_sc_hd__a21oi_1 _06716_ (.A1(_01687_),
    .A2(_01688_),
    .B1(net107),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _06717_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net77),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _06718_ (.A(net1044),
    .B(_01632_),
    .Y(_01690_));
 sky130_fd_sc_hd__a21oi_1 _06719_ (.A1(_01689_),
    .A2(_01690_),
    .B1(net105),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _06720_ (.A(net1257),
    .B(_01632_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01628_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand3b_1 _06722_ (.A_N(net103),
    .B(_01691_),
    .C(_01692_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_01628_),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(net212),
    .B(_01632_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21oi_1 _06725_ (.A1(_01693_),
    .A2(_01694_),
    .B1(net104),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _06726_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01628_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _06727_ (.A(net427),
    .B(_01632_),
    .Y(_01696_));
 sky130_fd_sc_hd__a21oi_1 _06728_ (.A1(_01695_),
    .A2(_01696_),
    .B1(net105),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _06729_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net77),
    .Y(_01697_));
 sky130_fd_sc_hd__nand2_1 _06730_ (.A(net705),
    .B(_01632_),
    .Y(_01698_));
 sky130_fd_sc_hd__a21oi_1 _06731_ (.A1(_01697_),
    .A2(_01698_),
    .B1(net107),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _06732_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_01628_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(net319),
    .B(_01632_),
    .Y(_01700_));
 sky130_fd_sc_hd__a21oi_1 _06734_ (.A1(_01699_),
    .A2(_01700_),
    .B1(net103),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01628_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _06736_ (.A(net932),
    .B(_01632_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21oi_1 _06737_ (.A1(_01701_),
    .A2(_01702_),
    .B1(net103),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _06738_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net77),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(net988),
    .B(_01632_),
    .Y(_01704_));
 sky130_fd_sc_hd__a21oi_1 _06740_ (.A1(_01703_),
    .A2(_01704_),
    .B1(net103),
    .Y(_00191_));
 sky130_fd_sc_hd__nor2_8 _06741_ (.A(_01396_),
    .B(_01474_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_8 _06742_ (.A(_01174_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_515 ();
 sky130_fd_sc_hd__nand2_1 _06744_ (.A(net1204),
    .B(_01706_),
    .Y(_01708_));
 sky130_fd_sc_hd__nor3_4 _06745_ (.A(_01162_),
    .B(_01396_),
    .C(_01474_),
    .Y(_01709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_514 ();
 sky130_fd_sc_hd__nand2_1 _06747_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net75),
    .Y(_01711_));
 sky130_fd_sc_hd__nand3b_1 _06748_ (.A_N(net104),
    .B(_01708_),
    .C(_01711_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net74),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _06750_ (.A(net731),
    .B(_01706_),
    .Y(_01713_));
 sky130_fd_sc_hd__a21oi_1 _06751_ (.A1(_01712_),
    .A2(_01713_),
    .B1(net105),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _06752_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net74),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _06753_ (.A(net305),
    .B(_01706_),
    .Y(_01715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_512 ();
 sky130_fd_sc_hd__a21oi_1 _06756_ (.A1(_01714_),
    .A2(_01715_),
    .B1(CPU_reset_a4),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _06757_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net75),
    .Y(_01718_));
 sky130_fd_sc_hd__nand2_1 _06758_ (.A(net828),
    .B(_01706_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_1 _06759_ (.A1(_01718_),
    .A2(_01719_),
    .B1(net107),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net74),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _06761_ (.A(net413),
    .B(_01706_),
    .Y(_01721_));
 sky130_fd_sc_hd__a21oi_1 _06762_ (.A1(_01720_),
    .A2(_01721_),
    .B1(net107),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net75),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _06764_ (.A(net311),
    .B(_01706_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_1 _06765_ (.A1(_01722_),
    .A2(_01723_),
    .B1(net106),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _06766_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net74),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_1 _06767_ (.A(net1028),
    .B(_01706_),
    .Y(_01725_));
 sky130_fd_sc_hd__a21oi_1 _06768_ (.A1(_01724_),
    .A2(_01725_),
    .B1(net104),
    .Y(_00198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_511 ();
 sky130_fd_sc_hd__nand2_1 _06770_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(_01709_),
    .Y(_01727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_510 ();
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(net1210),
    .B(_01706_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_1 _06773_ (.A1(_01727_),
    .A2(_01729_),
    .B1(net105),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net75),
    .Y(_01730_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(net1125),
    .B(_01706_),
    .Y(_01731_));
 sky130_fd_sc_hd__a21oi_1 _06776_ (.A1(_01730_),
    .A2(_01731_),
    .B1(net102),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net75),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _06778_ (.A(net1099),
    .B(_01706_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _06779_ (.A1(_01732_),
    .A2(_01733_),
    .B1(net106),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net74),
    .Y(_01734_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(net375),
    .B(_01706_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21oi_1 _06782_ (.A1(_01734_),
    .A2(_01735_),
    .B1(net106),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(net1136),
    .B(_01706_),
    .Y(_01736_));
 sky130_fd_sc_hd__nand2_1 _06784_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01709_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand3b_1 _06785_ (.A_N(net103),
    .B(_01736_),
    .C(_01737_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net75),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _06787_ (.A(net405),
    .B(_01706_),
    .Y(_01739_));
 sky130_fd_sc_hd__a21oi_1 _06788_ (.A1(_01738_),
    .A2(_01739_),
    .B1(net102),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _06789_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(_01709_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _06790_ (.A(net982),
    .B(_01706_),
    .Y(_01741_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_509 ();
 sky130_fd_sc_hd__a21oi_1 _06792_ (.A1(_01740_),
    .A2(_01741_),
    .B1(net104),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net74),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _06794_ (.A(net874),
    .B(_01706_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21oi_1 _06795_ (.A1(_01743_),
    .A2(_01744_),
    .B1(CPU_reset_a4),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _06796_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net75),
    .Y(_01745_));
 sky130_fd_sc_hd__nand2_1 _06797_ (.A(net1024),
    .B(_01706_),
    .Y(_01746_));
 sky130_fd_sc_hd__a21oi_1 _06798_ (.A1(_01745_),
    .A2(_01746_),
    .B1(net104),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _06799_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net74),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _06800_ (.A(net293),
    .B(_01706_),
    .Y(_01748_));
 sky130_fd_sc_hd__a21oi_1 _06801_ (.A1(_01747_),
    .A2(_01748_),
    .B1(CPU_reset_a4),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net74),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _06803_ (.A(net872),
    .B(_01706_),
    .Y(_01750_));
 sky130_fd_sc_hd__a21oi_1 _06804_ (.A1(_01749_),
    .A2(_01750_),
    .B1(net106),
    .Y(_00209_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_508 ();
 sky130_fd_sc_hd__nand2_1 _06806_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net74),
    .Y(_01752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_507 ();
 sky130_fd_sc_hd__nand2_1 _06808_ (.A(net660),
    .B(_01706_),
    .Y(_01754_));
 sky130_fd_sc_hd__a21oi_1 _06809_ (.A1(_01752_),
    .A2(_01754_),
    .B1(CPU_reset_a4),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net74),
    .Y(_01755_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(net425),
    .B(_01706_),
    .Y(_01756_));
 sky130_fd_sc_hd__a21oi_1 _06812_ (.A1(_01755_),
    .A2(_01756_),
    .B1(net105),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _06813_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net74),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(net217),
    .B(_01706_),
    .Y(_01758_));
 sky130_fd_sc_hd__a21oi_1 _06815_ (.A1(_01757_),
    .A2(_01758_),
    .B1(net102),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _06816_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net75),
    .Y(_01759_));
 sky130_fd_sc_hd__nand2_1 _06817_ (.A(net970),
    .B(_01706_),
    .Y(_01760_));
 sky130_fd_sc_hd__a21oi_1 _06818_ (.A1(_01759_),
    .A2(_01760_),
    .B1(net107),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _06819_ (.A(net1316),
    .B(_01706_),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01709_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand3b_1 _06821_ (.A_N(net103),
    .B(_01761_),
    .C(_01762_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _06822_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net74),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(net858),
    .B(_01706_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21oi_1 _06824_ (.A1(_01763_),
    .A2(_01764_),
    .B1(net107),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _06825_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net74),
    .Y(_01765_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(net1132),
    .B(_01706_),
    .Y(_01766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_506 ();
 sky130_fd_sc_hd__a21oi_1 _06828_ (.A1(_01765_),
    .A2(_01766_),
    .B1(net105),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(net1053),
    .B(_01706_),
    .Y(_01768_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01709_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand3b_1 _06831_ (.A_N(net103),
    .B(_01768_),
    .C(_01769_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net75),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _06833_ (.A(net509),
    .B(_01706_),
    .Y(_01771_));
 sky130_fd_sc_hd__a21oi_1 _06834_ (.A1(_01770_),
    .A2(_01771_),
    .B1(net104),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01709_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _06836_ (.A(net954),
    .B(_01706_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21oi_1 _06837_ (.A1(_01772_),
    .A2(_01773_),
    .B1(net103),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net74),
    .Y(_01774_));
 sky130_fd_sc_hd__nand2_1 _06839_ (.A(net1143),
    .B(_01706_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_1 _06840_ (.A1(_01774_),
    .A2(_01775_),
    .B1(CPU_reset_a4),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net75),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_1 _06842_ (.A(net721),
    .B(_01706_),
    .Y(_01777_));
 sky130_fd_sc_hd__a21oi_1 _06843_ (.A1(_01776_),
    .A2(_01777_),
    .B1(net104),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _06844_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01709_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(net725),
    .B(_01706_),
    .Y(_01779_));
 sky130_fd_sc_hd__a21oi_1 _06846_ (.A1(_01778_),
    .A2(_01779_),
    .B1(net103),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _06847_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_01709_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _06848_ (.A(net803),
    .B(_01706_),
    .Y(_01781_));
 sky130_fd_sc_hd__a21oi_1 _06849_ (.A1(_01780_),
    .A2(_01781_),
    .B1(net103),
    .Y(_00223_));
 sky130_fd_sc_hd__nor3_4 _06850_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01551_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_8 _06851_ (.A(_01174_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_505 ();
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(net1114),
    .B(_01783_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor4_4 _06854_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01162_),
    .D(_01551_),
    .Y(_01786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_504 ();
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net71),
    .Y(_01788_));
 sky130_fd_sc_hd__nand3b_1 _06857_ (.A_N(net104),
    .B(_01785_),
    .C(_01788_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net69),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _06859_ (.A(net612),
    .B(_01783_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21oi_1 _06860_ (.A1(_01789_),
    .A2(_01790_),
    .B1(net107),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net69),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(net926),
    .B(_01783_),
    .Y(_01792_));
 sky130_fd_sc_hd__a21oi_1 _06863_ (.A1(_01791_),
    .A2(_01792_),
    .B1(CPU_reset_a4),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net70),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(net757),
    .B(_01783_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21oi_1 _06866_ (.A1(_01793_),
    .A2(_01794_),
    .B1(net107),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net70),
    .Y(_01795_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(net223),
    .B(_01783_),
    .Y(_01796_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_503 ();
 sky130_fd_sc_hd__a21oi_1 _06870_ (.A1(_01795_),
    .A2(_01796_),
    .B1(net106),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _06871_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net70),
    .Y(_01798_));
 sky130_fd_sc_hd__nand2_1 _06872_ (.A(net261),
    .B(_01783_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21oi_1 _06873_ (.A1(_01798_),
    .A2(_01799_),
    .B1(net106),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _06874_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net69),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _06875_ (.A(net733),
    .B(_01783_),
    .Y(_01801_));
 sky130_fd_sc_hd__a21oi_1 _06876_ (.A1(_01800_),
    .A2(_01801_),
    .B1(net105),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net71),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(net391),
    .B(_01783_),
    .Y(_01803_));
 sky130_fd_sc_hd__a21oi_1 _06879_ (.A1(_01802_),
    .A2(_01803_),
    .B1(net104),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net70),
    .Y(_01804_));
 sky130_fd_sc_hd__nand2_1 _06881_ (.A(net571),
    .B(_01783_),
    .Y(_01805_));
 sky130_fd_sc_hd__a21oi_1 _06882_ (.A1(_01804_),
    .A2(_01805_),
    .B1(net102),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _06883_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net70),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _06884_ (.A(net373),
    .B(_01783_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21oi_1 _06885_ (.A1(_01806_),
    .A2(_01807_),
    .B1(net106),
    .Y(_00233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_502 ();
 sky130_fd_sc_hd__nand2_1 _06887_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net70),
    .Y(_01809_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_501 ();
 sky130_fd_sc_hd__nand2_1 _06889_ (.A(net1187),
    .B(_01783_),
    .Y(_01811_));
 sky130_fd_sc_hd__a21oi_1 _06890_ (.A1(_01809_),
    .A2(_01811_),
    .B1(net106),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01786_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(net882),
    .B(_01783_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21oi_1 _06893_ (.A1(_01812_),
    .A2(_01813_),
    .B1(net103),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net70),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_1 _06895_ (.A(net928),
    .B(_01783_),
    .Y(_01815_));
 sky130_fd_sc_hd__a21oi_1 _06896_ (.A1(_01814_),
    .A2(_01815_),
    .B1(net102),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _06897_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net71),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(net799),
    .B(_01783_),
    .Y(_01817_));
 sky130_fd_sc_hd__a21oi_1 _06899_ (.A1(_01816_),
    .A2(_01817_),
    .B1(net104),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net71),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(net1000),
    .B(_01783_),
    .Y(_01819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_500 ();
 sky130_fd_sc_hd__a21oi_1 _06903_ (.A1(_01818_),
    .A2(_01819_),
    .B1(net106),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net70),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _06905_ (.A(net1085),
    .B(_01783_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21oi_1 _06906_ (.A1(_01821_),
    .A2(_01822_),
    .B1(net102),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _06907_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net70),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _06908_ (.A(net549),
    .B(_01783_),
    .Y(_01824_));
 sky130_fd_sc_hd__a21oi_1 _06909_ (.A1(_01823_),
    .A2(_01824_),
    .B1(CPU_reset_a4),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net71),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _06911_ (.A(net597),
    .B(_01783_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21oi_1 _06912_ (.A1(_01825_),
    .A2(_01826_),
    .B1(net106),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _06913_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net69),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _06914_ (.A(net610),
    .B(_01783_),
    .Y(_01828_));
 sky130_fd_sc_hd__a21oi_1 _06915_ (.A1(_01827_),
    .A2(_01828_),
    .B1(CPU_reset_a4),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _06916_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net69),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _06917_ (.A(net389),
    .B(_01783_),
    .Y(_01830_));
 sky130_fd_sc_hd__a21oi_1 _06918_ (.A1(_01829_),
    .A2(_01830_),
    .B1(net105),
    .Y(_00243_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_499 ();
 sky130_fd_sc_hd__nand2_1 _06920_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net71),
    .Y(_01832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_498 ();
 sky130_fd_sc_hd__nand2_1 _06922_ (.A(net938),
    .B(_01783_),
    .Y(_01834_));
 sky130_fd_sc_hd__a21oi_1 _06923_ (.A1(_01832_),
    .A2(_01834_),
    .B1(net107),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _06924_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net71),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(net698),
    .B(_01783_),
    .Y(_01836_));
 sky130_fd_sc_hd__a21oi_1 _06926_ (.A1(_01835_),
    .A2(_01836_),
    .B1(net107),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _06927_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01786_),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _06928_ (.A(net690),
    .B(_01783_),
    .Y(_01838_));
 sky130_fd_sc_hd__a21oi_1 _06929_ (.A1(_01837_),
    .A2(_01838_),
    .B1(net103),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _06930_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net69),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(net644),
    .B(_01783_),
    .Y(_01840_));
 sky130_fd_sc_hd__a21oi_1 _06932_ (.A1(_01839_),
    .A2(_01840_),
    .B1(net107),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net69),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _06934_ (.A(net297),
    .B(_01783_),
    .Y(_01842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_497 ();
 sky130_fd_sc_hd__a21oi_1 _06936_ (.A1(_01841_),
    .A2(_01842_),
    .B1(net105),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _06937_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01786_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _06938_ (.A(net565),
    .B(_01783_),
    .Y(_01845_));
 sky130_fd_sc_hd__a21oi_1 _06939_ (.A1(_01844_),
    .A2(_01845_),
    .B1(net103),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _06940_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net70),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _06941_ (.A(net561),
    .B(_01783_),
    .Y(_01847_));
 sky130_fd_sc_hd__a21oi_1 _06942_ (.A1(_01846_),
    .A2(_01847_),
    .B1(net104),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01786_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _06944_ (.A(net958),
    .B(_01783_),
    .Y(_01849_));
 sky130_fd_sc_hd__a21oi_1 _06945_ (.A1(_01848_),
    .A2(_01849_),
    .B1(net105),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _06946_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net69),
    .Y(_01850_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(net976),
    .B(_01783_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21oi_1 _06948_ (.A1(_01850_),
    .A2(_01851_),
    .B1(net107),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _06949_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net70),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _06950_ (.A(net868),
    .B(_01783_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21oi_1 _06951_ (.A1(_01852_),
    .A2(_01853_),
    .B1(net104),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _06952_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01786_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _06953_ (.A(net525),
    .B(_01783_),
    .Y(_01855_));
 sky130_fd_sc_hd__a21oi_1 _06954_ (.A1(_01854_),
    .A2(_01855_),
    .B1(net103),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _06955_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_01786_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(net707),
    .B(_01783_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21oi_1 _06957_ (.A1(_01856_),
    .A2(_01857_),
    .B1(net103),
    .Y(_00255_));
 sky130_fd_sc_hd__nor4_4 _06958_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01162_),
    .D(_01315_),
    .Y(_01858_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_496 ();
 sky130_fd_sc_hd__nand2_1 _06960_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net67),
    .Y(_01860_));
 sky130_fd_sc_hd__nor3_4 _06961_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01315_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand2_8 _06962_ (.A(_01174_),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_495 ();
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(net715),
    .B(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21oi_1 _06965_ (.A1(_01860_),
    .A2(_01864_),
    .B1(net104),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net66),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(net924),
    .B(_01862_),
    .Y(_01866_));
 sky130_fd_sc_hd__a21oi_1 _06968_ (.A1(_01865_),
    .A2(_01866_),
    .B1(net105),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net66),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(net767),
    .B(_01862_),
    .Y(_01868_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_494 ();
 sky130_fd_sc_hd__a21oi_1 _06972_ (.A1(_01867_),
    .A2(_01868_),
    .B1(net106),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _06973_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net67),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _06974_ (.A(net793),
    .B(_01862_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21oi_1 _06975_ (.A1(_01870_),
    .A2(_01871_),
    .B1(net107),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net66),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _06977_ (.A(net986),
    .B(_01862_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21oi_1 _06978_ (.A1(_01872_),
    .A2(_01873_),
    .B1(net107),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _06979_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net67),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _06980_ (.A(net692),
    .B(_01862_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_1 _06981_ (.A1(_01874_),
    .A2(_01875_),
    .B1(net107),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _06982_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net67),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _06983_ (.A(net817),
    .B(_01862_),
    .Y(_01877_));
 sky130_fd_sc_hd__a21oi_1 _06984_ (.A1(_01876_),
    .A2(_01877_),
    .B1(net102),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net68),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _06986_ (.A(net395),
    .B(_01862_),
    .Y(_01879_));
 sky130_fd_sc_hd__a21oi_1 _06987_ (.A1(_01878_),
    .A2(_01879_),
    .B1(net105),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _06988_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net67),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _06989_ (.A(net367),
    .B(_01862_),
    .Y(_01881_));
 sky130_fd_sc_hd__a21oi_1 _06990_ (.A1(_01880_),
    .A2(_01881_),
    .B1(net102),
    .Y(_00264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_493 ();
 sky130_fd_sc_hd__nand2_1 _06992_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net66),
    .Y(_01883_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_492 ();
 sky130_fd_sc_hd__nand2_1 _06994_ (.A(net735),
    .B(_01862_),
    .Y(_01885_));
 sky130_fd_sc_hd__a21oi_1 _06995_ (.A1(_01883_),
    .A2(_01885_),
    .B1(net106),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _06996_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net66),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _06997_ (.A(net1010),
    .B(_01862_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21oi_1 _06998_ (.A1(_01886_),
    .A2(_01887_),
    .B1(CPU_reset_a4),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _06999_ (.A(net1259),
    .B(_01862_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01858_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand3b_1 _07001_ (.A_N(net103),
    .B(_01888_),
    .C(_01889_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _07002_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net67),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(net303),
    .B(_01862_),
    .Y(_01891_));
 sky130_fd_sc_hd__a21oi_1 _07004_ (.A1(_01890_),
    .A2(_01891_),
    .B1(net102),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net67),
    .Y(_01892_));
 sky130_fd_sc_hd__nand2_1 _07006_ (.A(net577),
    .B(_01862_),
    .Y(_01893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_491 ();
 sky130_fd_sc_hd__a21oi_1 _07008_ (.A1(_01892_),
    .A2(_01893_),
    .B1(net104),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _07009_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net66),
    .Y(_01895_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(net974),
    .B(_01862_),
    .Y(_01896_));
 sky130_fd_sc_hd__a21oi_1 _07011_ (.A1(_01895_),
    .A2(_01896_),
    .B1(net106),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net67),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _07013_ (.A(net523),
    .B(_01862_),
    .Y(_01898_));
 sky130_fd_sc_hd__a21oi_1 _07014_ (.A1(_01897_),
    .A2(_01898_),
    .B1(net102),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _07015_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net66),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _07016_ (.A(net468),
    .B(_01862_),
    .Y(_01900_));
 sky130_fd_sc_hd__a21oi_1 _07017_ (.A1(_01899_),
    .A2(_01900_),
    .B1(net106),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _07018_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net66),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(net301),
    .B(_01862_),
    .Y(_01902_));
 sky130_fd_sc_hd__a21oi_1 _07020_ (.A1(_01901_),
    .A2(_01902_),
    .B1(net106),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _07021_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net66),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _07022_ (.A(net600),
    .B(_01862_),
    .Y(_01904_));
 sky130_fd_sc_hd__a21oi_1 _07023_ (.A1(_01903_),
    .A2(_01904_),
    .B1(net106),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net68),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _07025_ (.A(net397),
    .B(_01862_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21oi_1 _07026_ (.A1(_01905_),
    .A2(_01906_),
    .B1(net105),
    .Y(_00275_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_490 ();
 sky130_fd_sc_hd__nand2_1 _07028_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net68),
    .Y(_01908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_489 ();
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(net703),
    .B(_01862_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21oi_1 _07031_ (.A1(_01908_),
    .A2(_01910_),
    .B1(net104),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _07032_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net67),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _07033_ (.A(net962),
    .B(_01862_),
    .Y(_01912_));
 sky130_fd_sc_hd__a21oi_1 _07034_ (.A1(_01911_),
    .A2(_01912_),
    .B1(net107),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _07035_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01858_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(net1004),
    .B(_01862_),
    .Y(_01914_));
 sky130_fd_sc_hd__a21oi_1 _07037_ (.A1(_01913_),
    .A2(_01914_),
    .B1(net103),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _07038_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net66),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _07039_ (.A(net773),
    .B(_01862_),
    .Y(_01916_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_488 ();
 sky130_fd_sc_hd__a21oi_1 _07041_ (.A1(_01915_),
    .A2(_01916_),
    .B1(net107),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _07042_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net68),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_1 _07043_ (.A(net1026),
    .B(_01862_),
    .Y(_01919_));
 sky130_fd_sc_hd__a21oi_1 _07044_ (.A1(_01918_),
    .A2(_01919_),
    .B1(net105),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01858_),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_1 _07046_ (.A(net513),
    .B(_01862_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21oi_1 _07047_ (.A1(_01920_),
    .A2(_01921_),
    .B1(net103),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_01858_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(net484),
    .B(_01862_),
    .Y(_01923_));
 sky130_fd_sc_hd__a21oi_1 _07050_ (.A1(_01922_),
    .A2(_01923_),
    .B1(net104),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01858_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _07052_ (.A(net1199),
    .B(_01862_),
    .Y(_01925_));
 sky130_fd_sc_hd__a21oi_1 _07053_ (.A1(_01924_),
    .A2(_01925_),
    .B1(net105),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _07054_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net66),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _07055_ (.A(net755),
    .B(_01862_),
    .Y(_01927_));
 sky130_fd_sc_hd__a21oi_1 _07056_ (.A1(_01926_),
    .A2(_01927_),
    .B1(net106),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _07057_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net67),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _07058_ (.A(net854),
    .B(_01862_),
    .Y(_01929_));
 sky130_fd_sc_hd__a21oi_1 _07059_ (.A1(_01928_),
    .A2(_01929_),
    .B1(net104),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _07060_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01858_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(net279),
    .B(_01862_),
    .Y(_01931_));
 sky130_fd_sc_hd__a21oi_1 _07062_ (.A1(_01930_),
    .A2(_01931_),
    .B1(net103),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net68),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(net1154),
    .B(_01862_),
    .Y(_01933_));
 sky130_fd_sc_hd__a21oi_1 _07065_ (.A1(_01932_),
    .A2(_01933_),
    .B1(net105),
    .Y(_00287_));
 sky130_fd_sc_hd__nor3_4 _07066_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01396_),
    .Y(_01934_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_487 ();
 sky130_fd_sc_hd__nand2_8 _07068_ (.A(_01174_),
    .B(_01934_),
    .Y(_01936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_486 ();
 sky130_fd_sc_hd__nand2_1 _07070_ (.A(net1413),
    .B(_01936_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor4_4 _07071_ (.A(\CPU_dmem_addr_a4[2] ),
    .B(\CPU_dmem_addr_a4[3] ),
    .C(_01162_),
    .D(_01396_),
    .Y(_01939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_485 ();
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net59),
    .Y(_01941_));
 sky130_fd_sc_hd__nand3b_1 _07074_ (.A_N(net104),
    .B(_01938_),
    .C(_01941_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _07075_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net60),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _07076_ (.A(net273),
    .B(_01936_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21oi_1 _07077_ (.A1(_01942_),
    .A2(_01943_),
    .B1(net105),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _07078_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net60),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _07079_ (.A(net381),
    .B(_01936_),
    .Y(_01945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_484 ();
 sky130_fd_sc_hd__a21oi_1 _07081_ (.A1(_01944_),
    .A2(_01945_),
    .B1(net106),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _07082_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net59),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(net325),
    .B(_01936_),
    .Y(_01948_));
 sky130_fd_sc_hd__a21oi_1 _07084_ (.A1(_01947_),
    .A2(_01948_),
    .B1(net107),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _07085_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net59),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _07086_ (.A(net676),
    .B(_01936_),
    .Y(_01950_));
 sky130_fd_sc_hd__a21oi_1 _07087_ (.A1(_01949_),
    .A2(_01950_),
    .B1(net106),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _07088_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net60),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _07089_ (.A(net1038),
    .B(_01936_),
    .Y(_01952_));
 sky130_fd_sc_hd__a21oi_1 _07090_ (.A1(_01951_),
    .A2(_01952_),
    .B1(net107),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net61),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _07092_ (.A(net825),
    .B(_01936_),
    .Y(_01954_));
 sky130_fd_sc_hd__a21oi_1 _07093_ (.A1(_01953_),
    .A2(_01954_),
    .B1(net102),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _07094_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net61),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _07095_ (.A(net998),
    .B(_01936_),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_1 _07096_ (.A1(_01955_),
    .A2(_01956_),
    .B1(net105),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net59),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _07098_ (.A(net864),
    .B(_01936_),
    .Y(_01958_));
 sky130_fd_sc_hd__a21oi_1 _07099_ (.A1(_01957_),
    .A2(_01958_),
    .B1(net102),
    .Y(_00296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_483 ();
 sky130_fd_sc_hd__nand2_1 _07101_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net59),
    .Y(_01960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_482 ();
 sky130_fd_sc_hd__nand2_1 _07103_ (.A(net894),
    .B(_01936_),
    .Y(_01962_));
 sky130_fd_sc_hd__a21oi_1 _07104_ (.A1(_01960_),
    .A2(_01962_),
    .B1(net106),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _07105_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net60),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(net531),
    .B(_01936_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21oi_1 _07107_ (.A1(_01963_),
    .A2(_01964_),
    .B1(CPU_reset_a4),
    .Y(_00298_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_481 ();
 sky130_fd_sc_hd__nand2_1 _07109_ (.A(net1249),
    .B(_01936_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_01939_),
    .Y(_01967_));
 sky130_fd_sc_hd__nand3b_1 _07111_ (.A_N(net103),
    .B(_01966_),
    .C(_01967_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net59),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _07113_ (.A(net237),
    .B(_01936_),
    .Y(_01969_));
 sky130_fd_sc_hd__a21oi_1 _07114_ (.A1(_01968_),
    .A2(_01969_),
    .B1(net102),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net61),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(net277),
    .B(_01936_),
    .Y(_01971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_479 ();
 sky130_fd_sc_hd__a21oi_1 _07119_ (.A1(_01970_),
    .A2(_01971_),
    .B1(net104),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _07120_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net60),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _07121_ (.A(net1063),
    .B(_01936_),
    .Y(_01975_));
 sky130_fd_sc_hd__a21oi_1 _07122_ (.A1(_01974_),
    .A2(_01975_),
    .B1(net106),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _07123_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net59),
    .Y(_01976_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(net905),
    .B(_01936_),
    .Y(_01977_));
 sky130_fd_sc_hd__a21oi_1 _07125_ (.A1(_01976_),
    .A2(_01977_),
    .B1(net104),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net60),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(net231),
    .B(_01936_),
    .Y(_01979_));
 sky130_fd_sc_hd__a21oi_1 _07128_ (.A1(_01978_),
    .A2(_01979_),
    .B1(CPU_reset_a4),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _07129_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net59),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(net1020),
    .B(_01936_),
    .Y(_01981_));
 sky130_fd_sc_hd__a21oi_1 _07131_ (.A1(_01980_),
    .A2(_01981_),
    .B1(net106),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net60),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _07133_ (.A(net289),
    .B(_01936_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21oi_1 _07134_ (.A1(_01982_),
    .A2(_01983_),
    .B1(CPU_reset_a4),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _07135_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net60),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(net1067),
    .B(_01936_),
    .Y(_01985_));
 sky130_fd_sc_hd__a21oi_1 _07137_ (.A1(_01984_),
    .A2(_01985_),
    .B1(net105),
    .Y(_00307_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_478 ();
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net60),
    .Y(_01987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_477 ();
 sky130_fd_sc_hd__nand2_1 _07141_ (.A(net444),
    .B(_01936_),
    .Y(_01989_));
 sky130_fd_sc_hd__a21oi_1 _07142_ (.A1(_01987_),
    .A2(_01989_),
    .B1(net107),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net59),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _07144_ (.A(net243),
    .B(_01936_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21oi_1 _07145_ (.A1(_01990_),
    .A2(_01991_),
    .B1(net107),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _07146_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_01939_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand2_1 _07147_ (.A(net1107),
    .B(_01936_),
    .Y(_01993_));
 sky130_fd_sc_hd__a21oi_1 _07148_ (.A1(_01992_),
    .A2(_01993_),
    .B1(net103),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _07149_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net60),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(net944),
    .B(_01936_),
    .Y(_01995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_476 ();
 sky130_fd_sc_hd__a21oi_1 _07152_ (.A1(_01994_),
    .A2(_01995_),
    .B1(net107),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net61),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_1 _07154_ (.A(net1116),
    .B(_01936_),
    .Y(_01998_));
 sky130_fd_sc_hd__a21oi_1 _07155_ (.A1(_01997_),
    .A2(_01998_),
    .B1(net105),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_01939_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(net547),
    .B(_01936_),
    .Y(_02000_));
 sky130_fd_sc_hd__a21oi_1 _07158_ (.A1(_01999_),
    .A2(_02000_),
    .B1(net103),
    .Y(_00313_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net59),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _07160_ (.A(net327),
    .B(_01936_),
    .Y(_02002_));
 sky130_fd_sc_hd__a21oi_1 _07161_ (.A1(_02001_),
    .A2(_02002_),
    .B1(net104),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _07162_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_01939_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _07163_ (.A(net860),
    .B(_01936_),
    .Y(_02004_));
 sky130_fd_sc_hd__a21oi_1 _07164_ (.A1(_02003_),
    .A2(_02004_),
    .B1(net105),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net60),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(net1164),
    .B(_01936_),
    .Y(_02006_));
 sky130_fd_sc_hd__a21oi_1 _07167_ (.A1(_02005_),
    .A2(_02006_),
    .B1(net106),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net59),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(net1119),
    .B(_01936_),
    .Y(_02008_));
 sky130_fd_sc_hd__a21oi_1 _07170_ (.A1(_02007_),
    .A2(_02008_),
    .B1(net104),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _07171_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_01939_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _07172_ (.A(net870),
    .B(_01936_),
    .Y(_02010_));
 sky130_fd_sc_hd__a21oi_1 _07173_ (.A1(_02009_),
    .A2(_02010_),
    .B1(net103),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _07174_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net61),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _07175_ (.A(net313),
    .B(_01936_),
    .Y(_02012_));
 sky130_fd_sc_hd__a21oi_1 _07176_ (.A1(_02011_),
    .A2(_02012_),
    .B1(net104),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2b_4 _07177_ (.A_N(\CPU_dmem_addr_a4[3] ),
    .B(\CPU_dmem_addr_a4[2] ),
    .Y(_02013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_475 ();
 sky130_fd_sc_hd__nor4_4 _07179_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_01162_),
    .D(_02013_),
    .Y(_02015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_474 ();
 sky130_fd_sc_hd__nand2_1 _07181_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(_02015_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor3_4 _07182_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_02013_),
    .Y(_02018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_473 ();
 sky130_fd_sc_hd__nand2_8 _07184_ (.A(_01174_),
    .B(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_472 ();
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(net1050),
    .B(_02020_),
    .Y(_02022_));
 sky130_fd_sc_hd__a21oi_1 _07187_ (.A1(_02017_),
    .A2(_02022_),
    .B1(net104),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _07188_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net57),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(net966),
    .B(_02020_),
    .Y(_02024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_471 ();
 sky130_fd_sc_hd__a21oi_1 _07191_ (.A1(_02023_),
    .A2(_02024_),
    .B1(net105),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _07192_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net57),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _07193_ (.A(net878),
    .B(_02020_),
    .Y(_02027_));
 sky130_fd_sc_hd__a21oi_1 _07194_ (.A1(_02026_),
    .A2(_02027_),
    .B1(net106),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _07195_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net56),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(net1261),
    .B(_02020_),
    .Y(_02029_));
 sky130_fd_sc_hd__a21oi_1 _07197_ (.A1(_02028_),
    .A2(_02029_),
    .B1(net107),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _07198_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net56),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _07199_ (.A(net569),
    .B(_02020_),
    .Y(_02031_));
 sky130_fd_sc_hd__a21oi_1 _07200_ (.A1(_02030_),
    .A2(_02031_),
    .B1(net106),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _07201_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net56),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _07202_ (.A(net608),
    .B(_02020_),
    .Y(_02033_));
 sky130_fd_sc_hd__a21oi_1 _07203_ (.A1(_02032_),
    .A2(_02033_),
    .B1(net107),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _07204_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net57),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(net573),
    .B(_02020_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21oi_1 _07206_ (.A1(_02034_),
    .A2(_02035_),
    .B1(net102),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _07207_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(_02015_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(net423),
    .B(_02020_),
    .Y(_02037_));
 sky130_fd_sc_hd__a21oi_1 _07209_ (.A1(_02036_),
    .A2(_02037_),
    .B1(net105),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _07210_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net56),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(net333),
    .B(_02020_),
    .Y(_02039_));
 sky130_fd_sc_hd__a21oi_1 _07212_ (.A1(_02038_),
    .A2(_02039_),
    .B1(net102),
    .Y(_00328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_470 ();
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net56),
    .Y(_02041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_469 ();
 sky130_fd_sc_hd__nand2_1 _07216_ (.A(net719),
    .B(_02020_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _07217_ (.A1(_02041_),
    .A2(_02043_),
    .B1(net106),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _07218_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net56),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(net911),
    .B(_02020_),
    .Y(_02045_));
 sky130_fd_sc_hd__a21oi_1 _07220_ (.A1(_02044_),
    .A2(_02045_),
    .B1(CPU_reset_a4),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(net58),
    .Y(_02046_));
 sky130_fd_sc_hd__nand2_1 _07222_ (.A(net271),
    .B(_02020_),
    .Y(_02047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_468 ();
 sky130_fd_sc_hd__a21oi_1 _07224_ (.A1(_02046_),
    .A2(_02047_),
    .B1(net103),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _07225_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net56),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_1 _07226_ (.A(net888),
    .B(_02020_),
    .Y(_02050_));
 sky130_fd_sc_hd__a21oi_1 _07227_ (.A1(_02049_),
    .A2(_02050_),
    .B1(net102),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net57),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(net686),
    .B(_02020_),
    .Y(_02052_));
 sky130_fd_sc_hd__a21oi_1 _07230_ (.A1(_02051_),
    .A2(_02052_),
    .B1(net104),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _07231_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net57),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(net309),
    .B(_02020_),
    .Y(_02054_));
 sky130_fd_sc_hd__a21oi_1 _07233_ (.A1(_02053_),
    .A2(_02054_),
    .B1(CPU_reset_a4),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net56),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _07235_ (.A(net579),
    .B(_02020_),
    .Y(_02056_));
 sky130_fd_sc_hd__a21oi_1 _07236_ (.A1(_02055_),
    .A2(_02056_),
    .B1(net102),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _07237_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net56),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(net202),
    .B(_02020_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21oi_1 _07239_ (.A1(_02057_),
    .A2(_02058_),
    .B1(CPU_reset_a4),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _07240_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net56),
    .Y(_02059_));
 sky130_fd_sc_hd__nand2_1 _07241_ (.A(net960),
    .B(_02020_),
    .Y(_02060_));
 sky130_fd_sc_hd__a21oi_1 _07242_ (.A1(_02059_),
    .A2(_02060_),
    .B1(net106),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _07243_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net57),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(net281),
    .B(_02020_),
    .Y(_02062_));
 sky130_fd_sc_hd__a21oi_1 _07245_ (.A1(_02061_),
    .A2(_02062_),
    .B1(net106),
    .Y(_00338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_467 ();
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net57),
    .Y(_02064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_466 ();
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(net1254),
    .B(_02020_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21oi_1 _07250_ (.A1(_02064_),
    .A2(_02066_),
    .B1(net105),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _07251_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net57),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _07252_ (.A(net807),
    .B(_02020_),
    .Y(_02068_));
 sky130_fd_sc_hd__a21oi_1 _07253_ (.A1(_02067_),
    .A2(_02068_),
    .B1(net102),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net56),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _07255_ (.A(net496),
    .B(_02020_),
    .Y(_02070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_465 ();
 sky130_fd_sc_hd__a21oi_1 _07257_ (.A1(_02069_),
    .A2(_02070_),
    .B1(net107),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(net1071),
    .B(_02020_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(net58),
    .Y(_02073_));
 sky130_fd_sc_hd__nand3b_1 _07260_ (.A_N(net103),
    .B(_02072_),
    .C(_02073_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _07261_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net57),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(net263),
    .B(_02020_),
    .Y(_02075_));
 sky130_fd_sc_hd__a21oi_1 _07263_ (.A1(_02074_),
    .A2(_02075_),
    .B1(net107),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(_02015_),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(net1069),
    .B(_02020_),
    .Y(_02077_));
 sky130_fd_sc_hd__a21oi_1 _07266_ (.A1(_02076_),
    .A2(_02077_),
    .B1(net105),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(net58),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(net830),
    .B(_02020_),
    .Y(_02079_));
 sky130_fd_sc_hd__a21oi_1 _07269_ (.A1(_02078_),
    .A2(_02079_),
    .B1(net103),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _07270_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net58),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _07271_ (.A(net821),
    .B(_02020_),
    .Y(_02081_));
 sky130_fd_sc_hd__a21oi_1 _07272_ (.A1(_02080_),
    .A2(_02081_),
    .B1(net103),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _07273_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(net58),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(net1040),
    .B(_02020_),
    .Y(_02083_));
 sky130_fd_sc_hd__a21oi_1 _07275_ (.A1(_02082_),
    .A2(_02083_),
    .B1(net105),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _07276_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net57),
    .Y(_02084_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(net1158),
    .B(_02020_),
    .Y(_02085_));
 sky130_fd_sc_hd__a21oi_1 _07278_ (.A1(_02084_),
    .A2(_02085_),
    .B1(net107),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _07279_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net56),
    .Y(_02086_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(net759),
    .B(_02020_),
    .Y(_02087_));
 sky130_fd_sc_hd__a21oi_1 _07281_ (.A1(_02086_),
    .A2(_02087_),
    .B1(net104),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(net58),
    .Y(_02088_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(net486),
    .B(_02020_),
    .Y(_02089_));
 sky130_fd_sc_hd__a21oi_1 _07284_ (.A1(_02088_),
    .A2(_02089_),
    .B1(net103),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _07285_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_02015_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _07286_ (.A(net1362),
    .B(_02020_),
    .Y(_02091_));
 sky130_fd_sc_hd__a21oi_1 _07287_ (.A1(_02090_),
    .A2(_02091_),
    .B1(net103),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_8 _07288_ (.A(_01551_),
    .B(_02013_),
    .Y(_02092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_464 ();
 sky130_fd_sc_hd__nand2_8 _07290_ (.A(_01174_),
    .B(_02092_),
    .Y(_02094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_463 ();
 sky130_fd_sc_hd__nand2_1 _07292_ (.A(net1313),
    .B(_02094_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor3_4 _07293_ (.A(_01162_),
    .B(_01551_),
    .C(_02013_),
    .Y(_02097_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_462 ();
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net53),
    .Y(_02099_));
 sky130_fd_sc_hd__nand3b_1 _07296_ (.A_N(net104),
    .B(_02096_),
    .C(_02099_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _07297_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net52),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(net1310),
    .B(_02094_),
    .Y(_02101_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_461 ();
 sky130_fd_sc_hd__a21oi_1 _07300_ (.A1(_02100_),
    .A2(_02101_),
    .B1(net105),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _07301_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net52),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(net688),
    .B(_02094_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21oi_1 _07303_ (.A1(_02103_),
    .A2(_02104_),
    .B1(net106),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net53),
    .Y(_02105_));
 sky130_fd_sc_hd__nand2_1 _07305_ (.A(net593),
    .B(_02094_),
    .Y(_02106_));
 sky130_fd_sc_hd__a21oi_1 _07306_ (.A1(_02105_),
    .A2(_02106_),
    .B1(net107),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net53),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _07308_ (.A(net464),
    .B(_02094_),
    .Y(_02108_));
 sky130_fd_sc_hd__a21oi_1 _07309_ (.A1(_02107_),
    .A2(_02108_),
    .B1(net106),
    .Y(_00356_));
 sky130_fd_sc_hd__nand2_1 _07310_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net53),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _07311_ (.A(net1180),
    .B(_02094_),
    .Y(_02110_));
 sky130_fd_sc_hd__a21oi_1 _07312_ (.A1(_02109_),
    .A2(_02110_),
    .B1(net106),
    .Y(_00357_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net52),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _07314_ (.A(net353),
    .B(_02094_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21oi_1 _07315_ (.A1(_02111_),
    .A2(_02112_),
    .B1(net102),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(_02097_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _07317_ (.A(net709),
    .B(_02094_),
    .Y(_02114_));
 sky130_fd_sc_hd__a21oi_1 _07318_ (.A1(_02113_),
    .A2(_02114_),
    .B1(net105),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _07319_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net52),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(net604),
    .B(_02094_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21oi_1 _07321_ (.A1(_02115_),
    .A2(_02116_),
    .B1(net104),
    .Y(_00360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_460 ();
 sky130_fd_sc_hd__nand2_1 _07323_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net53),
    .Y(_02118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_459 ();
 sky130_fd_sc_hd__nand2_1 _07325_ (.A(net494),
    .B(_02094_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21oi_1 _07326_ (.A1(_02118_),
    .A2(_02120_),
    .B1(net106),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net52),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _07328_ (.A(net1036),
    .B(_02094_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21oi_1 _07329_ (.A1(_02121_),
    .A2(_02122_),
    .B1(net106),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _07330_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(net53),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _07331_ (.A(net934),
    .B(_02094_),
    .Y(_02124_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_458 ();
 sky130_fd_sc_hd__a21oi_1 _07333_ (.A1(_02123_),
    .A2(_02124_),
    .B1(net103),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _07334_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net53),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(net206),
    .B(_02094_),
    .Y(_02127_));
 sky130_fd_sc_hd__a21oi_1 _07336_ (.A1(_02126_),
    .A2(_02127_),
    .B1(net102),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _07337_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net52),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _07338_ (.A(net765),
    .B(_02094_),
    .Y(_02129_));
 sky130_fd_sc_hd__a21oi_1 _07339_ (.A1(_02128_),
    .A2(_02129_),
    .B1(net104),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net52),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _07341_ (.A(net462),
    .B(_02094_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21oi_1 _07342_ (.A1(_02130_),
    .A2(_02131_),
    .B1(net106),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net53),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _07344_ (.A(net723),
    .B(_02094_),
    .Y(_02133_));
 sky130_fd_sc_hd__a21oi_1 _07345_ (.A1(_02132_),
    .A2(_02133_),
    .B1(net102),
    .Y(_00367_));
 sky130_fd_sc_hd__nand2_1 _07346_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net52),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(net363),
    .B(_02094_),
    .Y(_02135_));
 sky130_fd_sc_hd__a21oi_1 _07348_ (.A1(_02134_),
    .A2(_02135_),
    .B1(net106),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net52),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(net797),
    .B(_02094_),
    .Y(_02137_));
 sky130_fd_sc_hd__a21oi_1 _07351_ (.A1(_02136_),
    .A2(_02137_),
    .B1(net106),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net52),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _07353_ (.A(net915),
    .B(_02094_),
    .Y(_02139_));
 sky130_fd_sc_hd__a21oi_1 _07354_ (.A1(_02138_),
    .A2(_02139_),
    .B1(net107),
    .Y(_00370_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_457 ();
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net52),
    .Y(_02141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_456 ();
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(net1273),
    .B(_02094_),
    .Y(_02143_));
 sky130_fd_sc_hd__a21oi_1 _07359_ (.A1(_02141_),
    .A2(_02143_),
    .B1(net105),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net52),
    .Y(_02144_));
 sky130_fd_sc_hd__nand2_1 _07361_ (.A(net433),
    .B(_02094_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21oi_1 _07362_ (.A1(_02144_),
    .A2(_02145_),
    .B1(net102),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_1 _07363_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net52),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _07364_ (.A(net1002),
    .B(_02094_),
    .Y(_02147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_455 ();
 sky130_fd_sc_hd__a21oi_1 _07366_ (.A1(_02146_),
    .A2(_02147_),
    .B1(net107),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _07367_ (.A(net1191),
    .B(_02094_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_02097_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand3b_1 _07369_ (.A_N(net103),
    .B(_02149_),
    .C(_02150_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _07370_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net52),
    .Y(_02151_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(net769),
    .B(_02094_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21oi_1 _07372_ (.A1(_02151_),
    .A2(_02152_),
    .B1(net105),
    .Y(_00375_));
 sky130_fd_sc_hd__nand2_1 _07373_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net52),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _07374_ (.A(net1006),
    .B(_02094_),
    .Y(_02154_));
 sky130_fd_sc_hd__a21oi_1 _07375_ (.A1(_02153_),
    .A2(_02154_),
    .B1(net105),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_02097_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _07377_ (.A(net490),
    .B(_02094_),
    .Y(_02156_));
 sky130_fd_sc_hd__a21oi_1 _07378_ (.A1(_02155_),
    .A2(_02156_),
    .B1(net103),
    .Y(_00377_));
 sky130_fd_sc_hd__nand2_1 _07379_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net53),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _07380_ (.A(net674),
    .B(_02094_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_1 _07381_ (.A1(_02157_),
    .A2(_02158_),
    .B1(net103),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _07382_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_02097_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _07383_ (.A(net1097),
    .B(_02094_),
    .Y(_02160_));
 sky130_fd_sc_hd__a21oi_1 _07384_ (.A1(_02159_),
    .A2(_02160_),
    .B1(net105),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _07385_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net52),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(net385),
    .B(_02094_),
    .Y(_02162_));
 sky130_fd_sc_hd__a21oi_1 _07387_ (.A1(_02161_),
    .A2(_02162_),
    .B1(net106),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2_1 _07388_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net53),
    .Y(_02163_));
 sky130_fd_sc_hd__nand2_1 _07389_ (.A(net652),
    .B(_02094_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _07390_ (.A1(_02163_),
    .A2(_02164_),
    .B1(net103),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(net53),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _07392_ (.A(net771),
    .B(_02094_),
    .Y(_02166_));
 sky130_fd_sc_hd__a21oi_1 _07393_ (.A1(_02165_),
    .A2(_02166_),
    .B1(net103),
    .Y(_00382_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net53),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(net1229),
    .B(_02094_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21oi_1 _07396_ (.A1(_02167_),
    .A2(_02168_),
    .B1(net103),
    .Y(_00383_));
 sky130_fd_sc_hd__nor3_4 _07397_ (.A(_01162_),
    .B(_01315_),
    .C(_02013_),
    .Y(_02169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_454 ();
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net51),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_8 _07400_ (.A(_01315_),
    .B(_02013_),
    .Y(_02172_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_453 ();
 sky130_fd_sc_hd__nand2_8 _07402_ (.A(_01174_),
    .B(_02172_),
    .Y(_02174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_452 ();
 sky130_fd_sc_hd__nand2_1 _07404_ (.A(net650),
    .B(_02174_),
    .Y(_02176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_451 ();
 sky130_fd_sc_hd__a21oi_1 _07406_ (.A1(_02171_),
    .A2(_02176_),
    .B1(net104),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _07407_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net50),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(net339),
    .B(_02174_),
    .Y(_02179_));
 sky130_fd_sc_hd__a21oi_1 _07409_ (.A1(_02178_),
    .A2(_02179_),
    .B1(net107),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _07410_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net50),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _07411_ (.A(net225),
    .B(_02174_),
    .Y(_02181_));
 sky130_fd_sc_hd__a21oi_1 _07412_ (.A1(_02180_),
    .A2(_02181_),
    .B1(net106),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _07413_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net51),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(net269),
    .B(_02174_),
    .Y(_02183_));
 sky130_fd_sc_hd__a21oi_1 _07415_ (.A1(_02182_),
    .A2(_02183_),
    .B1(net102),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _07416_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net50),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _07417_ (.A(net1095),
    .B(_02174_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21oi_1 _07418_ (.A1(_02184_),
    .A2(_02185_),
    .B1(net106),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _07419_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net50),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _07420_ (.A(net221),
    .B(_02174_),
    .Y(_02187_));
 sky130_fd_sc_hd__a21oi_1 _07421_ (.A1(_02186_),
    .A2(_02187_),
    .B1(net107),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _07422_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net51),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _07423_ (.A(net421),
    .B(_02174_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_1 _07424_ (.A1(_02188_),
    .A2(_02189_),
    .B1(net104),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _07425_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net51),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(net846),
    .B(_02174_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21oi_1 _07427_ (.A1(_02190_),
    .A2(_02191_),
    .B1(net105),
    .Y(_00391_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_450 ();
 sky130_fd_sc_hd__nand2_1 _07429_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(_02169_),
    .Y(_02193_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_449 ();
 sky130_fd_sc_hd__nand2_1 _07431_ (.A(net345),
    .B(_02174_),
    .Y(_02195_));
 sky130_fd_sc_hd__a21oi_1 _07432_ (.A1(_02193_),
    .A2(_02195_),
    .B1(net102),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _07433_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net51),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _07434_ (.A(net331),
    .B(_02174_),
    .Y(_02197_));
 sky130_fd_sc_hd__a21oi_1 _07435_ (.A1(_02196_),
    .A2(_02197_),
    .B1(net106),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _07436_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net51),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _07437_ (.A(net618),
    .B(_02174_),
    .Y(_02199_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_448 ();
 sky130_fd_sc_hd__a21oi_1 _07439_ (.A1(_02198_),
    .A2(_02199_),
    .B1(CPU_reset_a4),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _07440_ (.A(net1178),
    .B(_02174_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _07441_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_02169_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand3b_1 _07442_ (.A_N(net103),
    .B(_02201_),
    .C(_02202_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(_02169_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _07444_ (.A(net684),
    .B(_02174_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21oi_1 _07445_ (.A1(_02203_),
    .A2(_02204_),
    .B1(net102),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net51),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(net208),
    .B(_02174_),
    .Y(_02206_));
 sky130_fd_sc_hd__a21oi_1 _07448_ (.A1(_02205_),
    .A2(_02206_),
    .B1(net104),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _07449_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net50),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _07450_ (.A(net747),
    .B(_02174_),
    .Y(_02208_));
 sky130_fd_sc_hd__a21oi_1 _07451_ (.A1(_02207_),
    .A2(_02208_),
    .B1(net106),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _07452_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_02169_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(net1141),
    .B(_02174_),
    .Y(_02210_));
 sky130_fd_sc_hd__a21oi_1 _07454_ (.A1(_02209_),
    .A2(_02210_),
    .B1(net104),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _07455_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net51),
    .Y(_02211_));
 sky130_fd_sc_hd__nand2_1 _07456_ (.A(net285),
    .B(_02174_),
    .Y(_02212_));
 sky130_fd_sc_hd__a21oi_1 _07457_ (.A1(_02211_),
    .A2(_02212_),
    .B1(CPU_reset_a4),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _07458_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net51),
    .Y(_02213_));
 sky130_fd_sc_hd__nand2_1 _07459_ (.A(net359),
    .B(_02174_),
    .Y(_02214_));
 sky130_fd_sc_hd__a21oi_1 _07460_ (.A1(_02213_),
    .A2(_02214_),
    .B1(net106),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _07461_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net50),
    .Y(_02215_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(net668),
    .B(_02174_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21oi_1 _07463_ (.A1(_02215_),
    .A2(_02216_),
    .B1(net107),
    .Y(_00402_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_447 ();
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net50),
    .Y(_02218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_446 ();
 sky130_fd_sc_hd__nand2_1 _07467_ (.A(net862),
    .B(_02174_),
    .Y(_02220_));
 sky130_fd_sc_hd__a21oi_1 _07468_ (.A1(_02218_),
    .A2(_02220_),
    .B1(net105),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _07469_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net50),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(net415),
    .B(_02174_),
    .Y(_02222_));
 sky130_fd_sc_hd__a21oi_1 _07471_ (.A1(_02221_),
    .A2(_02222_),
    .B1(net104),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net51),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _07473_ (.A(net662),
    .B(_02174_),
    .Y(_02224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_444 ();
 sky130_fd_sc_hd__a21oi_1 _07476_ (.A1(_02223_),
    .A2(_02224_),
    .B1(net107),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _07477_ (.A(net1032),
    .B(_02174_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand2_1 _07478_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_02169_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand3b_1 _07479_ (.A_N(net103),
    .B(_02227_),
    .C(_02228_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _07480_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net50),
    .Y(_02229_));
 sky130_fd_sc_hd__nand2_1 _07481_ (.A(net727),
    .B(_02174_),
    .Y(_02230_));
 sky130_fd_sc_hd__a21oi_1 _07482_ (.A1(_02229_),
    .A2(_02230_),
    .B1(net107),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net50),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _07484_ (.A(net287),
    .B(_02174_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_1 _07485_ (.A1(_02231_),
    .A2(_02232_),
    .B1(net105),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _07486_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_02169_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand2_1 _07487_ (.A(net642),
    .B(_02174_),
    .Y(_02234_));
 sky130_fd_sc_hd__a21oi_1 _07488_ (.A1(_02233_),
    .A2(_02234_),
    .B1(net103),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _07489_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_02169_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(net235),
    .B(_02174_),
    .Y(_02236_));
 sky130_fd_sc_hd__a21oi_1 _07491_ (.A1(_02235_),
    .A2(_02236_),
    .B1(net104),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_02169_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _07493_ (.A(net956),
    .B(_02174_),
    .Y(_02238_));
 sky130_fd_sc_hd__a21oi_1 _07494_ (.A1(_02237_),
    .A2(_02238_),
    .B1(net105),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net50),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _07496_ (.A(net907),
    .B(_02174_),
    .Y(_02240_));
 sky130_fd_sc_hd__a21oi_1 _07497_ (.A1(_02239_),
    .A2(_02240_),
    .B1(net107),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_02169_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _07499_ (.A(net507),
    .B(_02174_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21oi_1 _07500_ (.A1(_02241_),
    .A2(_02242_),
    .B1(net104),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_02169_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(net842),
    .B(_02174_),
    .Y(_02244_));
 sky130_fd_sc_hd__a21oi_1 _07503_ (.A1(_02243_),
    .A2(_02244_),
    .B1(net103),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _07504_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_02169_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_1 _07505_ (.A(net1630),
    .B(_02174_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21oi_1 _07506_ (.A1(_02245_),
    .A2(_02246_),
    .B1(net103),
    .Y(_00415_));
 sky130_fd_sc_hd__nor2_8 _07507_ (.A(_01396_),
    .B(_02013_),
    .Y(_02247_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_443 ();
 sky130_fd_sc_hd__nand2_8 _07509_ (.A(_01174_),
    .B(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_442 ();
 sky130_fd_sc_hd__nand2_1 _07511_ (.A(net1237),
    .B(_02249_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor3_4 _07512_ (.A(_01162_),
    .B(_01396_),
    .C(_02013_),
    .Y(_02252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_441 ();
 sky130_fd_sc_hd__nand2_1 _07514_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net48),
    .Y(_02254_));
 sky130_fd_sc_hd__nand3b_1 _07515_ (.A_N(net104),
    .B(_02251_),
    .C(_02254_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net49),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(net666),
    .B(_02249_),
    .Y(_02256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_440 ();
 sky130_fd_sc_hd__a21oi_1 _07519_ (.A1(_02255_),
    .A2(_02256_),
    .B1(net105),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net49),
    .Y(_02258_));
 sky130_fd_sc_hd__nand2_1 _07521_ (.A(net323),
    .B(_02249_),
    .Y(_02259_));
 sky130_fd_sc_hd__a21oi_1 _07522_ (.A1(_02258_),
    .A2(_02259_),
    .B1(CPU_reset_a4),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _07523_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net48),
    .Y(_02260_));
 sky130_fd_sc_hd__nand2_1 _07524_ (.A(net840),
    .B(_02249_),
    .Y(_02261_));
 sky130_fd_sc_hd__a21oi_1 _07525_ (.A1(_02260_),
    .A2(_02261_),
    .B1(net102),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _07526_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net48),
    .Y(_02262_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(net295),
    .B(_02249_),
    .Y(_02263_));
 sky130_fd_sc_hd__a21oi_1 _07528_ (.A1(_02262_),
    .A2(_02263_),
    .B1(net106),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _07529_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net48),
    .Y(_02264_));
 sky130_fd_sc_hd__nand2_1 _07530_ (.A(net1065),
    .B(_02249_),
    .Y(_02265_));
 sky130_fd_sc_hd__a21oi_1 _07531_ (.A1(_02264_),
    .A2(_02265_),
    .B1(net106),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net48),
    .Y(_02266_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(net583),
    .B(_02249_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _07534_ (.A1(_02266_),
    .A2(_02267_),
    .B1(net102),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _07535_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net49),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(net717),
    .B(_02249_),
    .Y(_02269_));
 sky130_fd_sc_hd__a21oi_1 _07537_ (.A1(_02268_),
    .A2(_02269_),
    .B1(net105),
    .Y(_00423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_439 ();
 sky130_fd_sc_hd__nand2_1 _07539_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net48),
    .Y(_02271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_438 ();
 sky130_fd_sc_hd__nand2_1 _07541_ (.A(net622),
    .B(_02249_),
    .Y(_02273_));
 sky130_fd_sc_hd__a21oi_1 _07542_ (.A1(_02271_),
    .A2(_02273_),
    .B1(net102),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net48),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _07544_ (.A(net498),
    .B(_02249_),
    .Y(_02275_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(_02274_),
    .A2(_02275_),
    .B1(net106),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _07546_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net48),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(net1145),
    .B(_02249_),
    .Y(_02277_));
 sky130_fd_sc_hd__a21oi_1 _07548_ (.A1(_02276_),
    .A2(_02277_),
    .B1(CPU_reset_a4),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _07549_ (.A(net1171),
    .B(_02249_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _07550_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_02252_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand3b_1 _07551_ (.A_N(net103),
    .B(_02278_),
    .C(_02279_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _07552_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(_02252_),
    .Y(_02280_));
 sky130_fd_sc_hd__nand2_1 _07553_ (.A(net307),
    .B(_02249_),
    .Y(_02281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_437 ();
 sky130_fd_sc_hd__a21oi_1 _07555_ (.A1(_02280_),
    .A2(_02281_),
    .B1(net102),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _07556_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net48),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(net636),
    .B(_02249_),
    .Y(_02284_));
 sky130_fd_sc_hd__a21oi_1 _07558_ (.A1(_02283_),
    .A2(_02284_),
    .B1(net104),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _07559_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net49),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(net616),
    .B(_02249_),
    .Y(_02286_));
 sky130_fd_sc_hd__a21oi_1 _07561_ (.A1(_02285_),
    .A2(_02286_),
    .B1(net106),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _07562_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(_02252_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(net1081),
    .B(_02249_),
    .Y(_02288_));
 sky130_fd_sc_hd__a21oi_1 _07564_ (.A1(_02287_),
    .A2(_02288_),
    .B1(net104),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _07565_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net49),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(net581),
    .B(_02249_),
    .Y(_02290_));
 sky130_fd_sc_hd__a21oi_1 _07567_ (.A1(_02289_),
    .A2(_02290_),
    .B1(net106),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net48),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _07569_ (.A(net440),
    .B(_02249_),
    .Y(_02292_));
 sky130_fd_sc_hd__a21oi_1 _07570_ (.A1(_02291_),
    .A2(_02292_),
    .B1(net106),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net49),
    .Y(_02293_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(net511),
    .B(_02249_),
    .Y(_02294_));
 sky130_fd_sc_hd__a21oi_1 _07573_ (.A1(_02293_),
    .A2(_02294_),
    .B1(net106),
    .Y(_00434_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_436 ();
 sky130_fd_sc_hd__nand2_1 _07575_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net49),
    .Y(_02296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_435 ();
 sky130_fd_sc_hd__nand2_1 _07577_ (.A(net215),
    .B(_02249_),
    .Y(_02298_));
 sky130_fd_sc_hd__a21oi_1 _07578_ (.A1(_02296_),
    .A2(_02298_),
    .B1(net105),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _07579_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net48),
    .Y(_02299_));
 sky130_fd_sc_hd__nand2_1 _07580_ (.A(net648),
    .B(_02249_),
    .Y(_02300_));
 sky130_fd_sc_hd__a21oi_1 _07581_ (.A1(_02299_),
    .A2(_02300_),
    .B1(net102),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _07582_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net48),
    .Y(_02301_));
 sky130_fd_sc_hd__nand2_1 _07583_ (.A(net521),
    .B(_02249_),
    .Y(_02302_));
 sky130_fd_sc_hd__a21oi_1 _07584_ (.A1(_02301_),
    .A2(_02302_),
    .B1(net107),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(net1079),
    .B(_02249_),
    .Y(_02303_));
 sky130_fd_sc_hd__nand2_1 _07586_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_02252_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand3b_1 _07587_ (.A_N(net103),
    .B(_02303_),
    .C(_02304_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _07588_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net49),
    .Y(_02305_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(net1090),
    .B(_02249_),
    .Y(_02306_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_434 ();
 sky130_fd_sc_hd__a21oi_1 _07591_ (.A1(_02305_),
    .A2(_02306_),
    .B1(net105),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net49),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(net283),
    .B(_02249_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21oi_1 _07594_ (.A1(_02308_),
    .A2(_02309_),
    .B1(net105),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _07595_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_02252_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand2_1 _07596_ (.A(net749),
    .B(_02249_),
    .Y(_02311_));
 sky130_fd_sc_hd__a21oi_1 _07597_ (.A1(_02310_),
    .A2(_02311_),
    .B1(net103),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_02252_),
    .Y(_02312_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(net502),
    .B(_02249_),
    .Y(_02313_));
 sky130_fd_sc_hd__a21oi_1 _07600_ (.A1(_02312_),
    .A2(_02313_),
    .B1(net104),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _07601_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_02252_),
    .Y(_02314_));
 sky130_fd_sc_hd__nand2_1 _07602_ (.A(net591),
    .B(_02249_),
    .Y(_02315_));
 sky130_fd_sc_hd__a21oi_1 _07603_ (.A1(_02314_),
    .A2(_02315_),
    .B1(net105),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net49),
    .Y(_02316_));
 sky130_fd_sc_hd__nand2_1 _07605_ (.A(net1123),
    .B(_02249_),
    .Y(_02317_));
 sky130_fd_sc_hd__a21oi_1 _07606_ (.A1(_02316_),
    .A2(_02317_),
    .B1(net107),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _07607_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(_02252_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _07608_ (.A(net317),
    .B(_02249_),
    .Y(_02319_));
 sky130_fd_sc_hd__a21oi_1 _07609_ (.A1(_02318_),
    .A2(_02319_),
    .B1(net103),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_02252_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _07611_ (.A(net247),
    .B(_02249_),
    .Y(_02321_));
 sky130_fd_sc_hd__a21oi_1 _07612_ (.A1(_02320_),
    .A2(_02321_),
    .B1(net103),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(_02252_),
    .Y(_02322_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(net379),
    .B(_02249_),
    .Y(_02323_));
 sky130_fd_sc_hd__a21oi_1 _07615_ (.A1(_02322_),
    .A2(_02323_),
    .B1(net103),
    .Y(_00447_));
 sky130_fd_sc_hd__nor4_4 _07616_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_01162_),
    .D(_01317_),
    .Y(_02324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_433 ();
 sky130_fd_sc_hd__nand2_1 _07618_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net46),
    .Y(_02326_));
 sky130_fd_sc_hd__nor3_4 _07619_ (.A(\CPU_dmem_addr_a4[0] ),
    .B(\CPU_dmem_addr_a4[1] ),
    .C(_01317_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_8 _07620_ (.A(_01174_),
    .B(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_432 ();
 sky130_fd_sc_hd__nand2_1 _07622_ (.A(net401),
    .B(_02328_),
    .Y(_02330_));
 sky130_fd_sc_hd__a21oi_1 _07623_ (.A1(_02326_),
    .A2(_02330_),
    .B1(net104),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _07624_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net47),
    .Y(_02331_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(net990),
    .B(_02328_),
    .Y(_02332_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_431 ();
 sky130_fd_sc_hd__a21oi_1 _07627_ (.A1(_02331_),
    .A2(_02332_),
    .B1(net107),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _07628_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net45),
    .Y(_02334_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(net435),
    .B(_02328_),
    .Y(_02335_));
 sky130_fd_sc_hd__a21oi_1 _07630_ (.A1(_02334_),
    .A2(_02335_),
    .B1(CPU_reset_a4),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net46),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(net474),
    .B(_02328_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21oi_1 _07633_ (.A1(_02336_),
    .A2(_02337_),
    .B1(net107),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _07634_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net45),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _07635_ (.A(net739),
    .B(_02328_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21oi_1 _07636_ (.A1(_02338_),
    .A2(_02339_),
    .B1(net106),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _07637_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net46),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(net255),
    .B(_02328_),
    .Y(_02341_));
 sky130_fd_sc_hd__a21oi_1 _07639_ (.A1(_02340_),
    .A2(_02341_),
    .B1(net106),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _07640_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net47),
    .Y(_02342_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(net267),
    .B(_02328_),
    .Y(_02343_));
 sky130_fd_sc_hd__a21oi_1 _07642_ (.A1(_02342_),
    .A2(_02343_),
    .B1(net102),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _07643_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net47),
    .Y(_02344_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(net1055),
    .B(_02328_),
    .Y(_02345_));
 sky130_fd_sc_hd__a21oi_1 _07645_ (.A1(_02344_),
    .A2(_02345_),
    .B1(net105),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _07646_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net46),
    .Y(_02346_));
 sky130_fd_sc_hd__nand2_1 _07647_ (.A(net321),
    .B(_02328_),
    .Y(_02347_));
 sky130_fd_sc_hd__a21oi_1 _07648_ (.A1(_02346_),
    .A2(_02347_),
    .B1(net102),
    .Y(_00456_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_430 ();
 sky130_fd_sc_hd__nand2_1 _07650_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net45),
    .Y(_02349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_429 ();
 sky130_fd_sc_hd__nand2_1 _07652_ (.A(net595),
    .B(_02328_),
    .Y(_02351_));
 sky130_fd_sc_hd__a21oi_1 _07653_ (.A1(_02349_),
    .A2(_02351_),
    .B1(net106),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net45),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _07655_ (.A(net448),
    .B(_02328_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21oi_1 _07656_ (.A1(_02352_),
    .A2(_02353_),
    .B1(CPU_reset_a4),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _07657_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_02324_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _07658_ (.A(net233),
    .B(_02328_),
    .Y(_02355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_428 ();
 sky130_fd_sc_hd__a21oi_1 _07660_ (.A1(_02354_),
    .A2(_02355_),
    .B1(net103),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net46),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(net638),
    .B(_02328_),
    .Y(_02358_));
 sky130_fd_sc_hd__a21oi_1 _07663_ (.A1(_02357_),
    .A2(_02358_),
    .B1(net102),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _07664_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net47),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(net403),
    .B(_02328_),
    .Y(_02360_));
 sky130_fd_sc_hd__a21oi_1 _07666_ (.A1(_02359_),
    .A2(_02360_),
    .B1(net104),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _07667_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net45),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _07668_ (.A(net743),
    .B(_02328_),
    .Y(_02362_));
 sky130_fd_sc_hd__a21oi_1 _07669_ (.A1(_02361_),
    .A2(_02362_),
    .B1(CPU_reset_a4),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _07670_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net46),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _07671_ (.A(net918),
    .B(_02328_),
    .Y(_02364_));
 sky130_fd_sc_hd__a21oi_1 _07672_ (.A1(_02363_),
    .A2(_02364_),
    .B1(net104),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net45),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _07674_ (.A(net936),
    .B(_02328_),
    .Y(_02366_));
 sky130_fd_sc_hd__a21oi_1 _07675_ (.A1(_02365_),
    .A2(_02366_),
    .B1(CPU_reset_a4),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _07676_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net45),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(net265),
    .B(_02328_),
    .Y(_02368_));
 sky130_fd_sc_hd__a21oi_1 _07678_ (.A1(_02367_),
    .A2(_02368_),
    .B1(net106),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net45),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(net972),
    .B(_02328_),
    .Y(_02370_));
 sky130_fd_sc_hd__a21oi_1 _07681_ (.A1(_02369_),
    .A2(_02370_),
    .B1(net106),
    .Y(_00466_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_427 ();
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net47),
    .Y(_02372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_426 ();
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(net852),
    .B(_02328_),
    .Y(_02374_));
 sky130_fd_sc_hd__a21oi_1 _07686_ (.A1(_02372_),
    .A2(_02374_),
    .B1(net105),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net47),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_1 _07688_ (.A(net886),
    .B(_02328_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21oi_1 _07689_ (.A1(_02375_),
    .A2(_02376_),
    .B1(net104),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _07690_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net46),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(net259),
    .B(_02328_),
    .Y(_02378_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_425 ();
 sky130_fd_sc_hd__a21oi_1 _07693_ (.A1(_02377_),
    .A2(_02378_),
    .B1(net107),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_02324_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _07695_ (.A(net626),
    .B(_02328_),
    .Y(_02381_));
 sky130_fd_sc_hd__a21oi_1 _07696_ (.A1(_02380_),
    .A2(_02381_),
    .B1(net103),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net47),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_1 _07698_ (.A(net892),
    .B(_02328_),
    .Y(_02383_));
 sky130_fd_sc_hd__a21oi_1 _07699_ (.A1(_02382_),
    .A2(_02383_),
    .B1(net107),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _07700_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net47),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _07701_ (.A(net1156),
    .B(_02328_),
    .Y(_02385_));
 sky130_fd_sc_hd__a21oi_1 _07702_ (.A1(_02384_),
    .A2(_02385_),
    .B1(net105),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(net1160),
    .B(_02328_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _07704_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_02324_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand3b_1 _07705_ (.A_N(net103),
    .B(_02386_),
    .C(_02387_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(net46),
    .Y(_02388_));
 sky130_fd_sc_hd__nand2_1 _07707_ (.A(net337),
    .B(_02328_),
    .Y(_02389_));
 sky130_fd_sc_hd__a21oi_1 _07708_ (.A1(_02388_),
    .A2(_02389_),
    .B1(net103),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_02324_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _07710_ (.A(net1166),
    .B(_02328_),
    .Y(_02391_));
 sky130_fd_sc_hd__a21oi_1 _07711_ (.A1(_02390_),
    .A2(_02391_),
    .B1(net105),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net45),
    .Y(_02392_));
 sky130_fd_sc_hd__nand2_1 _07713_ (.A(net811),
    .B(_02328_),
    .Y(_02393_));
 sky130_fd_sc_hd__a21oi_1 _07714_ (.A1(_02392_),
    .A2(_02393_),
    .B1(CPU_reset_a4),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net46),
    .Y(_02394_));
 sky130_fd_sc_hd__nand2_1 _07716_ (.A(net587),
    .B(_02328_),
    .Y(_02395_));
 sky130_fd_sc_hd__a21oi_1 _07717_ (.A1(_02394_),
    .A2(_02395_),
    .B1(net104),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _07718_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_02324_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_1 _07719_ (.A(net763),
    .B(_02328_),
    .Y(_02397_));
 sky130_fd_sc_hd__a21oi_1 _07720_ (.A1(_02396_),
    .A2(_02397_),
    .B1(net103),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net46),
    .Y(_02398_));
 sky130_fd_sc_hd__nand2_1 _07722_ (.A(net470),
    .B(_02328_),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_1 _07723_ (.A1(_02398_),
    .A2(_02399_),
    .B1(net105),
    .Y(_00479_));
 sky130_fd_sc_hd__nor2_8 _07724_ (.A(_01317_),
    .B(_01551_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_8 _07725_ (.A(_01174_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_424 ();
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(net1139),
    .B(_02401_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor3_4 _07728_ (.A(_01162_),
    .B(_01317_),
    .C(_01551_),
    .Y(_02404_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_423 ();
 sky130_fd_sc_hd__nand2_1 _07730_ (.A(\CPU_dmem_wr_data_a4[0] ),
    .B(net41),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3b_1 _07731_ (.A_N(net104),
    .B(_02403_),
    .C(_02406_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(\CPU_dmem_wr_data_a4[10] ),
    .B(net42),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(net1195),
    .B(_02401_),
    .Y(_02408_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_422 ();
 sky130_fd_sc_hd__a21oi_1 _07735_ (.A1(_02407_),
    .A2(_02408_),
    .B1(net105),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(\CPU_dmem_wr_data_a4[11] ),
    .B(net42),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(net791),
    .B(_02401_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21oi_1 _07738_ (.A1(_02410_),
    .A2(_02411_),
    .B1(CPU_reset_a4),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(\CPU_dmem_wr_data_a4[12] ),
    .B(net41),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _07740_ (.A(net239),
    .B(_02401_),
    .Y(_02413_));
 sky130_fd_sc_hd__a21oi_1 _07741_ (.A1(_02412_),
    .A2(_02413_),
    .B1(net102),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _07742_ (.A(\CPU_dmem_wr_data_a4[13] ),
    .B(net41),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(net527),
    .B(_02401_),
    .Y(_02415_));
 sky130_fd_sc_hd__a21oi_1 _07744_ (.A1(_02414_),
    .A2(_02415_),
    .B1(net106),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(\CPU_dmem_wr_data_a4[14] ),
    .B(net41),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(net219),
    .B(_02401_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21oi_1 _07747_ (.A1(_02416_),
    .A2(_02417_),
    .B1(net107),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(\CPU_dmem_wr_data_a4[15] ),
    .B(net42),
    .Y(_02418_));
 sky130_fd_sc_hd__nand2_1 _07749_ (.A(net1048),
    .B(_02401_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21oi_1 _07750_ (.A1(_02418_),
    .A2(_02419_),
    .B1(net105),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _07751_ (.A(\CPU_dmem_wr_data_a4[16] ),
    .B(net41),
    .Y(_02420_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(net245),
    .B(_02401_),
    .Y(_02421_));
 sky130_fd_sc_hd__a21oi_1 _07753_ (.A1(_02420_),
    .A2(_02421_),
    .B1(net104),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(\CPU_dmem_wr_data_a4[17] ),
    .B(net41),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _07755_ (.A(net948),
    .B(_02401_),
    .Y(_02423_));
 sky130_fd_sc_hd__a21oi_1 _07756_ (.A1(_02422_),
    .A2(_02423_),
    .B1(net102),
    .Y(_00488_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_421 ();
 sky130_fd_sc_hd__nand2_1 _07758_ (.A(\CPU_dmem_wr_data_a4[18] ),
    .B(net41),
    .Y(_02425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_420 ();
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(net567),
    .B(_02401_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21oi_1 _07761_ (.A1(_02425_),
    .A2(_02427_),
    .B1(net106),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(\CPU_dmem_wr_data_a4[19] ),
    .B(net42),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_1 _07763_ (.A(net563),
    .B(_02401_),
    .Y(_02429_));
 sky130_fd_sc_hd__a21oi_1 _07764_ (.A1(_02428_),
    .A2(_02429_),
    .B1(CPU_reset_a4),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(\CPU_dmem_wr_data_a4[1] ),
    .B(_02404_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _07766_ (.A(net251),
    .B(_02401_),
    .Y(_02431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_419 ();
 sky130_fd_sc_hd__a21oi_1 _07768_ (.A1(_02430_),
    .A2(_02431_),
    .B1(net103),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(\CPU_dmem_wr_data_a4[20] ),
    .B(net41),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _07770_ (.A(net204),
    .B(_02401_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21oi_1 _07771_ (.A1(_02433_),
    .A2(_02434_),
    .B1(net102),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _07772_ (.A(\CPU_dmem_wr_data_a4[21] ),
    .B(net41),
    .Y(_02435_));
 sky130_fd_sc_hd__nand2_1 _07773_ (.A(net1042),
    .B(_02401_),
    .Y(_02436_));
 sky130_fd_sc_hd__a21oi_1 _07774_ (.A1(_02435_),
    .A2(_02436_),
    .B1(net104),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _07775_ (.A(\CPU_dmem_wr_data_a4[22] ),
    .B(net42),
    .Y(_02437_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(net930),
    .B(_02401_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21oi_1 _07777_ (.A1(_02437_),
    .A2(_02438_),
    .B1(CPU_reset_a4),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _07778_ (.A(\CPU_dmem_wr_data_a4[23] ),
    .B(net41),
    .Y(_02439_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(net417),
    .B(_02401_),
    .Y(_02440_));
 sky130_fd_sc_hd__a21oi_1 _07780_ (.A1(_02439_),
    .A2(_02440_),
    .B1(net104),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _07781_ (.A(\CPU_dmem_wr_data_a4[24] ),
    .B(net42),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _07782_ (.A(net640),
    .B(_02401_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21oi_1 _07783_ (.A1(_02441_),
    .A2(_02442_),
    .B1(CPU_reset_a4),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _07784_ (.A(\CPU_dmem_wr_data_a4[25] ),
    .B(net41),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(net545),
    .B(_02401_),
    .Y(_02444_));
 sky130_fd_sc_hd__a21oi_1 _07786_ (.A1(_02443_),
    .A2(_02444_),
    .B1(net106),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _07787_ (.A(\CPU_dmem_wr_data_a4[26] ),
    .B(net42),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _07788_ (.A(net429),
    .B(_02401_),
    .Y(_02446_));
 sky130_fd_sc_hd__a21oi_1 _07789_ (.A1(_02445_),
    .A2(_02446_),
    .B1(net106),
    .Y(_00498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_418 ();
 sky130_fd_sc_hd__nand2_1 _07791_ (.A(\CPU_dmem_wr_data_a4[27] ),
    .B(net42),
    .Y(_02448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_417 ();
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(net836),
    .B(_02401_),
    .Y(_02450_));
 sky130_fd_sc_hd__a21oi_1 _07794_ (.A1(_02448_),
    .A2(_02450_),
    .B1(net105),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _07795_ (.A(\CPU_dmem_wr_data_a4[28] ),
    .B(net42),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _07796_ (.A(net795),
    .B(_02401_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21oi_1 _07797_ (.A1(_02451_),
    .A2(_02452_),
    .B1(net107),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _07798_ (.A(\CPU_dmem_wr_data_a4[29] ),
    .B(net41),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(net377),
    .B(_02401_),
    .Y(_02454_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_416 ();
 sky130_fd_sc_hd__a21oi_1 _07801_ (.A1(_02453_),
    .A2(_02454_),
    .B1(net107),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(\CPU_dmem_wr_data_a4[2] ),
    .B(_02404_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(net1341),
    .B(_02401_),
    .Y(_02457_));
 sky130_fd_sc_hd__a21oi_1 _07804_ (.A1(_02456_),
    .A2(_02457_),
    .B1(net103),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(\CPU_dmem_wr_data_a4[30] ),
    .B(net42),
    .Y(_02458_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(net210),
    .B(_02401_),
    .Y(_02459_));
 sky130_fd_sc_hd__a21oi_1 _07807_ (.A1(_02458_),
    .A2(_02459_),
    .B1(net107),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(\CPU_dmem_wr_data_a4[31] ),
    .B(net42),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _07809_ (.A(net634),
    .B(_02401_),
    .Y(_02461_));
 sky130_fd_sc_hd__a21oi_1 _07810_ (.A1(_02460_),
    .A2(_02461_),
    .B1(net105),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _07811_ (.A(net1321),
    .B(_02401_),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(\CPU_dmem_wr_data_a4[3] ),
    .B(_02404_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand3b_1 _07813_ (.A_N(net103),
    .B(_02462_),
    .C(_02463_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(\CPU_dmem_wr_data_a4[4] ),
    .B(_02404_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(net419),
    .B(_02401_),
    .Y(_02465_));
 sky130_fd_sc_hd__a21oi_1 _07816_ (.A1(_02464_),
    .A2(_02465_),
    .B1(net103),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(\CPU_dmem_wr_data_a4[5] ),
    .B(_02404_),
    .Y(_02466_));
 sky130_fd_sc_hd__nand2_1 _07818_ (.A(net832),
    .B(_02401_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21oi_1 _07819_ (.A1(_02466_),
    .A2(_02467_),
    .B1(net103),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(\CPU_dmem_wr_data_a4[6] ),
    .B(net42),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _07821_ (.A(net898),
    .B(_02401_),
    .Y(_02469_));
 sky130_fd_sc_hd__a21oi_1 _07822_ (.A1(_02468_),
    .A2(_02469_),
    .B1(CPU_reset_a4),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(\CPU_dmem_wr_data_a4[7] ),
    .B(net41),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _07824_ (.A(net535),
    .B(_02401_),
    .Y(_02471_));
 sky130_fd_sc_hd__a21oi_1 _07825_ (.A1(_02470_),
    .A2(_02471_),
    .B1(net104),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(\CPU_dmem_wr_data_a4[8] ),
    .B(_02404_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(net658),
    .B(_02401_),
    .Y(_02473_));
 sky130_fd_sc_hd__a21oi_1 _07828_ (.A1(_02472_),
    .A2(_02473_),
    .B1(net103),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(\CPU_dmem_wr_data_a4[9] ),
    .B(net41),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(net1352),
    .B(_02401_),
    .Y(_02475_));
 sky130_fd_sc_hd__a21oi_1 _07831_ (.A1(_02474_),
    .A2(_02475_),
    .B1(net105),
    .Y(_00511_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_414 ();
 sky130_fd_sc_hd__nor2b_1 _07834_ (.A(net108),
    .B_N(net1679),
    .Y(_00512_));
 sky130_fd_sc_hd__nor2b_1 _07835_ (.A(net108),
    .B_N(net1292),
    .Y(_00513_));
 sky130_fd_sc_hd__nor2b_1 _07836_ (.A(net109),
    .B_N(net1504),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2b_1 _07837_ (.A(CPU_reset_a3),
    .B_N(net1684),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2b_1 _07838_ (.A(net109),
    .B_N(net1503),
    .Y(_00516_));
 sky130_fd_sc_hd__nor2b_1 _07839_ (.A(net108),
    .B_N(net1269),
    .Y(_00517_));
 sky130_fd_sc_hd__nor2b_1 _07840_ (.A(net108),
    .B_N(net1307),
    .Y(_00518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_412 ();
 sky130_fd_sc_hd__nor2b_1 _07843_ (.A(net108),
    .B_N(net1312),
    .Y(_00519_));
 sky130_fd_sc_hd__nor2b_1 _07844_ (.A(net108),
    .B_N(net1418),
    .Y(_00520_));
 sky130_fd_sc_hd__nor2b_1 _07845_ (.A(net109),
    .B_N(net1610),
    .Y(_00521_));
 sky130_fd_sc_hd__nor2b_1 _07846_ (.A(net108),
    .B_N(net1409),
    .Y(_00522_));
 sky130_fd_sc_hd__nor2b_1 _07847_ (.A(CPU_reset_a3),
    .B_N(net1676),
    .Y(_00523_));
 sky130_fd_sc_hd__nor2b_1 _07848_ (.A(CPU_reset_a3),
    .B_N(net1675),
    .Y(_00524_));
 sky130_fd_sc_hd__nor2b_1 _07849_ (.A(net110),
    .B_N(net1671),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2b_1 _07850_ (.A(net108),
    .B_N(net1607),
    .Y(_00526_));
 sky130_fd_sc_hd__nor2b_1 _07851_ (.A(net110),
    .B_N(net1511),
    .Y(_00527_));
 sky130_fd_sc_hd__nor2b_1 _07852_ (.A(net109),
    .B_N(net1542),
    .Y(_00528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_411 ();
 sky130_fd_sc_hd__nor2b_1 _07854_ (.A(net108),
    .B_N(net1279),
    .Y(_00529_));
 sky130_fd_sc_hd__nor2b_1 _07855_ (.A(net109),
    .B_N(net1571),
    .Y(_00530_));
 sky130_fd_sc_hd__nor2b_1 _07856_ (.A(net110),
    .B_N(net1669),
    .Y(_00531_));
 sky130_fd_sc_hd__nor2b_1 _07857_ (.A(net108),
    .B_N(net1455),
    .Y(_00532_));
 sky130_fd_sc_hd__nor2b_1 _07858_ (.A(net108),
    .B_N(net1266),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2b_1 _07859_ (.A(CPU_reset_a3),
    .B_N(net1666),
    .Y(_00534_));
 sky130_fd_sc_hd__nor2b_1 _07860_ (.A(net109),
    .B_N(net1690),
    .Y(_00535_));
 sky130_fd_sc_hd__nor2b_1 _07861_ (.A(CPU_reset_a3),
    .B_N(net1683),
    .Y(_00536_));
 sky130_fd_sc_hd__nor2b_1 _07862_ (.A(CPU_reset_a3),
    .B_N(net1520),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2b_1 _07863_ (.A(net110),
    .B_N(net1673),
    .Y(_00538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_410 ();
 sky130_fd_sc_hd__nor2b_1 _07865_ (.A(CPU_reset_a3),
    .B_N(net1618),
    .Y(_00539_));
 sky130_fd_sc_hd__nor2b_1 _07866_ (.A(net110),
    .B_N(net1685),
    .Y(_00540_));
 sky130_fd_sc_hd__nor2b_1 _07867_ (.A(CPU_reset_a3),
    .B_N(net1689),
    .Y(_00541_));
 sky130_fd_sc_hd__nor2b_1 _07868_ (.A(CPU_reset_a3),
    .B_N(net1674),
    .Y(_00542_));
 sky130_fd_sc_hd__nor2b_1 _07869_ (.A(CPU_reset_a3),
    .B_N(net1678),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2b_1 _07870_ (.A_N(CPU_is_addi_a3),
    .B(CPU_is_slt_a3),
    .Y(_02482_));
 sky130_fd_sc_hd__nor2b_4 _07871_ (.A(CPU_is_addi_a3),
    .B_N(CPU_is_add_a3),
    .Y(_02483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_409 ();
 sky130_fd_sc_hd__a221oi_4 _07873_ (.A1(_05629_),
    .A2(_02482_),
    .B1(_02483_),
    .B2(_05636_),
    .C1(CPU_is_slti_a3),
    .Y(_02485_));
 sky130_fd_sc_hd__o21ai_1 _07874_ (.A1(_05525_),
    .A2(_05523_),
    .B1(CPU_is_slt_a3),
    .Y(_02486_));
 sky130_fd_sc_hd__nand4_1 _07875_ (.A(_05525_),
    .B(_01106_),
    .C(_01109_),
    .D(_02485_),
    .Y(_02487_));
 sky130_fd_sc_hd__a21oi_1 _07876_ (.A1(_01052_),
    .A2(_01102_),
    .B1(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _07877_ (.A(CPU_is_add_a3),
    .B(CPU_is_addi_a3),
    .Y(_02489_));
 sky130_fd_sc_hd__o21ai_2 _07878_ (.A1(_05523_),
    .A2(_05633_),
    .B1(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_407 ();
 sky130_fd_sc_hd__nand4_2 _07881_ (.A(_05633_),
    .B(_05567_),
    .C(_05572_),
    .D(_05800_),
    .Y(_02493_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_404 ();
 sky130_fd_sc_hd__nand4_1 _07885_ (.A(_05576_),
    .B(_05581_),
    .C(_05586_),
    .D(_05783_),
    .Y(_02497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_403 ();
 sky130_fd_sc_hd__inv_1 _07887_ (.A(_05739_),
    .Y(_02499_));
 sky130_fd_sc_hd__a21oi_1 _07888_ (.A1(_05599_),
    .A2(_05603_),
    .B1(_05598_),
    .Y(_02500_));
 sky130_fd_sc_hd__o21bai_1 _07889_ (.A1(_02499_),
    .A2(_02500_),
    .B1_N(_05738_),
    .Y(_02501_));
 sky130_fd_sc_hd__a21oi_1 _07890_ (.A1(_05594_),
    .A2(_02501_),
    .B1(_05593_),
    .Y(_02502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_400 ();
 sky130_fd_sc_hd__nand4_1 _07894_ (.A(_05590_),
    .B(_05748_),
    .C(_05757_),
    .D(_05766_),
    .Y(_02506_));
 sky130_fd_sc_hd__a21o_1 _07895_ (.A1(_05567_),
    .A2(_05571_),
    .B1(_05566_),
    .X(_02507_));
 sky130_fd_sc_hd__a21o_1 _07896_ (.A1(_05800_),
    .A2(_02507_),
    .B1(_05799_),
    .X(_02508_));
 sky130_fd_sc_hd__a21oi_1 _07897_ (.A1(_05633_),
    .A2(_02508_),
    .B1(_05632_),
    .Y(_02509_));
 sky130_fd_sc_hd__o41ai_1 _07898_ (.A1(_02493_),
    .A2(_02497_),
    .A3(_02502_),
    .A4(_02506_),
    .B1(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__or2_0 _07899_ (.A(_02493_),
    .B(_02497_),
    .X(_02511_));
 sky130_fd_sc_hd__inv_1 _07900_ (.A(_05766_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21oi_1 _07901_ (.A1(_05747_),
    .A2(_05757_),
    .B1(_05756_),
    .Y(_02513_));
 sky130_fd_sc_hd__o21bai_1 _07902_ (.A1(_02512_),
    .A2(_02513_),
    .B1_N(_05765_),
    .Y(_02514_));
 sky130_fd_sc_hd__a21oi_1 _07903_ (.A1(_05590_),
    .A2(_02514_),
    .B1(_05589_),
    .Y(_02515_));
 sky130_fd_sc_hd__inv_1 _07904_ (.A(_05783_),
    .Y(_02516_));
 sky130_fd_sc_hd__a21oi_1 _07905_ (.A1(_05581_),
    .A2(_05585_),
    .B1(_05580_),
    .Y(_02517_));
 sky130_fd_sc_hd__o21bai_1 _07906_ (.A1(_02516_),
    .A2(_02517_),
    .B1_N(_05782_),
    .Y(_02518_));
 sky130_fd_sc_hd__a21oi_1 _07907_ (.A1(_05576_),
    .A2(_02518_),
    .B1(_05575_),
    .Y(_02519_));
 sky130_fd_sc_hd__o22ai_1 _07908_ (.A1(_02511_),
    .A2(_02515_),
    .B1(_02519_),
    .B2(_02493_),
    .Y(_02520_));
 sky130_fd_sc_hd__nor3_2 _07909_ (.A(_02490_),
    .B(_02510_),
    .C(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__inv_1 _07910_ (.A(_05686_),
    .Y(_02522_));
 sky130_fd_sc_hd__clkinvlp_4 _07911_ (.A(_05695_),
    .Y(_02523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_398 ();
 sky130_fd_sc_hd__nand4_1 _07914_ (.A(_05608_),
    .B(_05704_),
    .C(_05713_),
    .D(_05722_),
    .Y(_02526_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(_05612_),
    .B(_05677_),
    .Y(_02527_));
 sky130_fd_sc_hd__or4_2 _07916_ (.A(_02522_),
    .B(_02523_),
    .C(_02526_),
    .D(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__inv_1 _07917_ (.A(_05668_),
    .Y(_02529_));
 sky130_fd_sc_hd__a21oi_1 _07918_ (.A1(_05649_),
    .A2(_05659_),
    .B1(_05658_),
    .Y(_02530_));
 sky130_fd_sc_hd__o21bai_1 _07919_ (.A1(_02529_),
    .A2(_02530_),
    .B1_N(_05667_),
    .Y(_02531_));
 sky130_fd_sc_hd__a21oi_1 _07920_ (.A1(_05616_),
    .A2(_02531_),
    .B1(_05615_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _07921_ (.A(_02528_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__inv_1 _07922_ (.A(_05619_),
    .Y(_02534_));
 sky130_fd_sc_hd__nor2b_1 _07923_ (.A(_05628_),
    .B_N(_05624_),
    .Y(_02535_));
 sky130_fd_sc_hd__o21a_1 _07924_ (.A1(_05623_),
    .A2(_02535_),
    .B1(_05641_),
    .X(_02536_));
 sky130_fd_sc_hd__o21ai_1 _07925_ (.A1(_05640_),
    .A2(_02536_),
    .B1(_05620_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand4_1 _07926_ (.A(_05616_),
    .B(_05650_),
    .C(_05659_),
    .D(_05668_),
    .Y(_02538_));
 sky130_fd_sc_hd__a211oi_1 _07927_ (.A1(_02534_),
    .A2(_02537_),
    .B1(_02538_),
    .C1(_02528_),
    .Y(_02539_));
 sky130_fd_sc_hd__a21oi_1 _07928_ (.A1(_05676_),
    .A2(_05686_),
    .B1(_05685_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21bai_1 _07929_ (.A1(_02523_),
    .A2(_02540_),
    .B1_N(_05694_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21oi_1 _07930_ (.A1(_05612_),
    .A2(_02541_),
    .B1(_05611_),
    .Y(_02542_));
 sky130_fd_sc_hd__clkinvlp_4 _07931_ (.A(_05722_),
    .Y(_02543_));
 sky130_fd_sc_hd__a21oi_1 _07932_ (.A1(_05703_),
    .A2(_05713_),
    .B1(_05712_),
    .Y(_02544_));
 sky130_fd_sc_hd__o21bai_1 _07933_ (.A1(_02543_),
    .A2(_02544_),
    .B1_N(_05721_),
    .Y(_02545_));
 sky130_fd_sc_hd__a21oi_1 _07934_ (.A1(_05608_),
    .A2(_02545_),
    .B1(_05607_),
    .Y(_02546_));
 sky130_fd_sc_hd__o21ai_0 _07935_ (.A1(_02526_),
    .A2(_02542_),
    .B1(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__nand4_1 _07936_ (.A(_05594_),
    .B(_05599_),
    .C(_05604_),
    .D(_05739_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor3_2 _07937_ (.A(_02511_),
    .B(_02506_),
    .C(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__o31ai_1 _07938_ (.A1(_02533_),
    .A2(_02539_),
    .A3(_02547_),
    .B1(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__inv_1 _07939_ (.A(CPU_is_slti_a3),
    .Y(_02551_));
 sky130_fd_sc_hd__mux2i_1 _07940_ (.A0(_02551_),
    .A1(_05636_),
    .S(CPU_is_add_a3),
    .Y(_02552_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(_05629_),
    .B(CPU_is_addi_a3),
    .Y(_02553_));
 sky130_fd_sc_hd__o21ai_1 _07942_ (.A1(CPU_is_addi_a3),
    .A2(_02552_),
    .B1(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand4_1 _07943_ (.A(_05620_),
    .B(_05624_),
    .C(_05629_),
    .D(_05641_),
    .Y(_02555_));
 sky130_fd_sc_hd__nor3_1 _07944_ (.A(_02528_),
    .B(_02538_),
    .C(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _07945_ (.A(_02549_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__a21oi_1 _07946_ (.A1(_05633_),
    .A2(_02557_),
    .B1(_02490_),
    .Y(_02558_));
 sky130_fd_sc_hd__a211oi_2 _07947_ (.A1(_02521_),
    .A2(_02550_),
    .B1(_02554_),
    .C1(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__a211oi_4 _07948_ (.A1(_02485_),
    .A2(_02486_),
    .B1(_02488_),
    .C1(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_397 ();
 sky130_fd_sc_hd__nand2b_1 _07950_ (.A_N(\CPU_rd_a5[2] ),
    .B(\CPU_rd_a5[3] ),
    .Y(_02562_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_396 ();
 sky130_fd_sc_hd__inv_1 _07952_ (.A(\CPU_rd_a3[2] ),
    .Y(_02564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_395 ();
 sky130_fd_sc_hd__nand3_2 _07954_ (.A(_02564_),
    .B(\CPU_rd_a3[3] ),
    .C(_01036_),
    .Y(_02566_));
 sky130_fd_sc_hd__o21a_4 _07955_ (.A1(_01036_),
    .A2(_02562_),
    .B1(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__clkinv_2 _07956_ (.A(CPU_valid_load_a5),
    .Y(_02568_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_394 ();
 sky130_fd_sc_hd__nor2_1 _07958_ (.A(\CPU_rd_a3[0] ),
    .B(\CPU_rd_a3[1] ),
    .Y(_02570_));
 sky130_fd_sc_hd__nor2_1 _07959_ (.A(\CPU_rd_a3[2] ),
    .B(\CPU_rd_a3[3] ),
    .Y(_02571_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(_02570_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__o211ai_4 _07961_ (.A1(\CPU_rd_a3[4] ),
    .A2(_02572_),
    .B1(_01036_),
    .C1(CPU_rd_valid_a3),
    .Y(_02573_));
 sky130_fd_sc_hd__o22ai_4 _07962_ (.A1(_02568_),
    .A2(\CPU_rd_a5[4] ),
    .B1(\CPU_rd_a3[4] ),
    .B2(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__nand2b_1 _07963_ (.A_N(\CPU_rd_a5[0] ),
    .B(\CPU_rd_a5[1] ),
    .Y(_02575_));
 sky130_fd_sc_hd__inv_1 _07964_ (.A(\CPU_rd_a3[0] ),
    .Y(_02576_));
 sky130_fd_sc_hd__nand3_1 _07965_ (.A(_02576_),
    .B(\CPU_rd_a3[1] ),
    .C(_01036_),
    .Y(_02577_));
 sky130_fd_sc_hd__o21ai_4 _07966_ (.A1(_01036_),
    .A2(_02575_),
    .B1(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_4 _07967_ (.A(_02574_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__nor2_8 _07968_ (.A(_02567_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__nor2_8 _07969_ (.A(CPU_reset_a3),
    .B(_01035_),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_8 _07970_ (.A(_02580_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_391 ();
 sky130_fd_sc_hd__clkinv_16 _07974_ (.A(net109),
    .Y(_02586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_390 ();
 sky130_fd_sc_hd__and3_2 _07976_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[0] ),
    .C(_01035_),
    .X(_02588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_387 ();
 sky130_fd_sc_hd__o21ai_4 _07980_ (.A1(_01036_),
    .A2(_02562_),
    .B1(_02566_),
    .Y(_02592_));
 sky130_fd_sc_hd__o22a_4 _07981_ (.A1(_02568_),
    .A2(\CPU_rd_a5[4] ),
    .B1(\CPU_rd_a3[4] ),
    .B2(_02573_),
    .X(_02593_));
 sky130_fd_sc_hd__o21a_2 _07982_ (.A1(_01036_),
    .A2(_02575_),
    .B1(_02577_),
    .X(_02594_));
 sky130_fd_sc_hd__nor2_8 _07983_ (.A(_02593_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_8 _07984_ (.A(_02592_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_386 ();
 sky130_fd_sc_hd__and3_1 _07986_ (.A(net1820),
    .B(net97),
    .C(_02596_),
    .X(_02598_));
 sky130_fd_sc_hd__a21oi_1 _07987_ (.A1(_02580_),
    .A2(_02588_),
    .B1(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__o21ai_0 _07988_ (.A1(_02560_),
    .A2(_02582_),
    .B1(_02599_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor3_2 _07989_ (.A(CPU_is_slti_a3),
    .B(CPU_is_slt_a3),
    .C(CPU_is_add_a3),
    .Y(_02600_));
 sky130_fd_sc_hd__nor2_8 _07990_ (.A(CPU_is_addi_a3),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_385 ();
 sky130_fd_sc_hd__nor2_2 _07992_ (.A(_05616_),
    .B(_05677_),
    .Y(_02603_));
 sky130_fd_sc_hd__nor3_2 _07993_ (.A(_05620_),
    .B(_05641_),
    .C(_05513_),
    .Y(_02604_));
 sky130_fd_sc_hd__nor2b_2 _07994_ (.A(_05620_),
    .B_N(_05642_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor3_2 _07995_ (.A(_05621_),
    .B(_02604_),
    .C(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nor2b_1 _07996_ (.A(_05659_),
    .B_N(_05651_),
    .Y(_02607_));
 sky130_fd_sc_hd__nor2_1 _07997_ (.A(_05660_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__o31ai_4 _07998_ (.A1(_05650_),
    .A2(_05659_),
    .A3(_02606_),
    .B1(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__nor2b_1 _07999_ (.A(_05686_),
    .B_N(_05678_),
    .Y(_02610_));
 sky130_fd_sc_hd__nor2_1 _08000_ (.A(_05687_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__nor2b_1 _08001_ (.A(_05616_),
    .B_N(_05669_),
    .Y(_02612_));
 sky130_fd_sc_hd__inv_1 _08002_ (.A(_05677_),
    .Y(_02613_));
 sky130_fd_sc_hd__o211ai_2 _08003_ (.A1(_05617_),
    .A2(_02612_),
    .B1(_02522_),
    .C1(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand2_1 _08004_ (.A(_02611_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__a41oi_1 _08005_ (.A1(_02529_),
    .A2(_02522_),
    .A3(_02603_),
    .A4(_02609_),
    .B1(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__xnor2_1 _08006_ (.A(_05695_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__a21oi_4 _08007_ (.A1(_01080_),
    .A2(_05673_),
    .B1(_05554_),
    .Y(_02618_));
 sky130_fd_sc_hd__inv_1 _08008_ (.A(_05690_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21oi_2 _08009_ (.A1(_05682_),
    .A2(_02619_),
    .B1(_05691_),
    .Y(_02620_));
 sky130_fd_sc_hd__o31ai_4 _08010_ (.A1(_05681_),
    .A2(_05690_),
    .A3(_02618_),
    .B1(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__o21ba_1 _08011_ (.A1(_05517_),
    .A2(_05645_),
    .B1_N(_05646_),
    .X(_02622_));
 sky130_fd_sc_hd__or4_4 _08012_ (.A(_05558_),
    .B(_05654_),
    .C(_05663_),
    .D(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__inv_1 _08013_ (.A(_05663_),
    .Y(_02624_));
 sky130_fd_sc_hd__nor2b_2 _08014_ (.A(_05654_),
    .B_N(_05559_),
    .Y(_02625_));
 sky130_fd_sc_hd__nor2b_1 _08015_ (.A(_05663_),
    .B_N(_05655_),
    .Y(_02626_));
 sky130_fd_sc_hd__a211oi_4 _08016_ (.A1(_02624_),
    .A2(_02625_),
    .B1(_02626_),
    .C1(_05664_),
    .Y(_02627_));
 sky130_fd_sc_hd__or3_2 _08017_ (.A(_05553_),
    .B(_05672_),
    .C(_05681_),
    .X(_02628_));
 sky130_fd_sc_hd__a211oi_4 _08018_ (.A1(_02623_),
    .A2(_02627_),
    .B1(_02628_),
    .C1(_05690_),
    .Y(_02629_));
 sky130_fd_sc_hd__or2_2 _08019_ (.A(_02621_),
    .B(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__xor2_2 _08020_ (.A(_05699_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__nand2b_4 _08021_ (.A_N(CPU_is_addi_a3),
    .B(CPU_is_add_a3),
    .Y(_02632_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_383 ();
 sky130_fd_sc_hd__o22ai_4 _08024_ (.A1(_02601_),
    .A2(_02617_),
    .B1(_02631_),
    .B2(_02632_),
    .Y(_02635_));
 sky130_fd_sc_hd__mux2_8 _08025_ (.A0(\CPU_dmem_rd_data_a5[10] ),
    .A1(_02635_),
    .S(_01036_),
    .X(_02636_));
 sky130_fd_sc_hd__nand2_1 _08026_ (.A(_02580_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_382 ();
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(net1356),
    .B(_02596_),
    .Y(_02639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__a21oi_1 _08030_ (.A1(_02637_),
    .A2(_02639_),
    .B1(net108),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(net1320),
    .B(_02596_),
    .Y(_02641_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__inv_1 _08034_ (.A(_05691_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_1 _08035_ (.A1(_05690_),
    .A2(_02644_),
    .B1(_05699_),
    .Y(_02645_));
 sky130_fd_sc_hd__nor2_2 _08036_ (.A(_05700_),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__nor2b_1 _08037_ (.A(_05562_),
    .B_N(_05637_),
    .Y(_02647_));
 sky130_fd_sc_hd__nor3_1 _08038_ (.A(_05558_),
    .B(_05645_),
    .C(_05654_),
    .Y(_02648_));
 sky130_fd_sc_hd__o21ai_2 _08039_ (.A1(_05563_),
    .A2(_02647_),
    .B1(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__nor3b_1 _08040_ (.A(_05558_),
    .B(_05654_),
    .C_N(_05646_),
    .Y(_02650_));
 sky130_fd_sc_hd__nor3_2 _08041_ (.A(_05655_),
    .B(_02625_),
    .C(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__a211oi_4 _08042_ (.A1(_02649_),
    .A2(_02651_),
    .B1(_05663_),
    .C1(_02628_),
    .Y(_02652_));
 sky130_fd_sc_hd__inv_1 _08043_ (.A(_05672_),
    .Y(_02653_));
 sky130_fd_sc_hd__a21oi_1 _08044_ (.A1(_05664_),
    .A2(_02653_),
    .B1(_05673_),
    .Y(_02654_));
 sky130_fd_sc_hd__inv_1 _08045_ (.A(_05681_),
    .Y(_02655_));
 sky130_fd_sc_hd__a21oi_1 _08046_ (.A1(_05554_),
    .A2(_02655_),
    .B1(_05682_),
    .Y(_02656_));
 sky130_fd_sc_hd__o31ai_4 _08047_ (.A1(_05553_),
    .A2(_05681_),
    .A3(_02654_),
    .B1(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__nor4_4 _08048_ (.A(_05691_),
    .B(_05700_),
    .C(_02652_),
    .D(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__or3_1 _08049_ (.A(_05548_),
    .B(_02646_),
    .C(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__o21ai_1 _08050_ (.A1(_02646_),
    .A2(_02658_),
    .B1(_05548_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand3_4 _08051_ (.A(_02483_),
    .B(_02659_),
    .C(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__a21oi_4 _08052_ (.A1(_05687_),
    .A2(_02523_),
    .B1(_05696_),
    .Y(_02662_));
 sky130_fd_sc_hd__a21o_1 _08053_ (.A1(_05617_),
    .A2(_02613_),
    .B1(_05678_),
    .X(_02663_));
 sky130_fd_sc_hd__nor2b_1 _08054_ (.A(_05668_),
    .B_N(_05660_),
    .Y(_02664_));
 sky130_fd_sc_hd__nor2_1 _08055_ (.A(_05669_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__inv_1 _08056_ (.A(_05650_),
    .Y(_02666_));
 sky130_fd_sc_hd__nor2b_1 _08057_ (.A(_05624_),
    .B_N(_05630_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2b_1 _08058_ (.A_N(_05642_),
    .B(_05641_),
    .Y(_02668_));
 sky130_fd_sc_hd__inv_1 _08059_ (.A(_05620_),
    .Y(_02669_));
 sky130_fd_sc_hd__o311a_1 _08060_ (.A1(_05625_),
    .A2(_05642_),
    .A3(_02667_),
    .B1(_02668_),
    .C1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__or2_0 _08061_ (.A(_05621_),
    .B(_05651_),
    .X(_02671_));
 sky130_fd_sc_hd__nor2_2 _08062_ (.A(_05659_),
    .B(_05668_),
    .Y(_02672_));
 sky130_fd_sc_hd__o221ai_4 _08063_ (.A1(_02666_),
    .A2(_05651_),
    .B1(_02670_),
    .B2(_02671_),
    .C1(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__a21boi_1 _08064_ (.A1(_02665_),
    .A2(_02673_),
    .B1_N(_02603_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand2_1 _08065_ (.A(_02522_),
    .B(_02523_),
    .Y(_02675_));
 sky130_fd_sc_hd__o21bai_2 _08066_ (.A1(_02663_),
    .A2(_02674_),
    .B1_N(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__clkinvlp_4 _08067_ (.A(_05612_),
    .Y(_02677_));
 sky130_fd_sc_hd__a211o_4 _08068_ (.A1(_02662_),
    .A2(_02676_),
    .B1(_02677_),
    .C1(_02601_),
    .X(_02678_));
 sky130_fd_sc_hd__or2_4 _08069_ (.A(CPU_is_addi_a3),
    .B(_02600_),
    .X(_02679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__nand4_4 _08071_ (.A(_02677_),
    .B(_02679_),
    .C(_02662_),
    .D(_02676_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_1 _08072_ (.A(\CPU_dmem_rd_data_a5[11] ),
    .B(_01036_),
    .Y(_02682_));
 sky130_fd_sc_hd__a41oi_4 _08073_ (.A1(_01036_),
    .A2(_02661_),
    .A3(_02678_),
    .A4(_02681_),
    .B1(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _08074_ (.A(_02580_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21oi_1 _08075_ (.A1(_02641_),
    .A2(_02684_),
    .B1(net109),
    .Y(_00546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__nand2b_1 _08078_ (.A_N(_05617_),
    .B(_05616_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor4_1 _08079_ (.A(_05612_),
    .B(_05677_),
    .C(_05686_),
    .D(_05695_),
    .Y(_02688_));
 sky130_fd_sc_hd__inv_1 _08080_ (.A(_05669_),
    .Y(_02689_));
 sky130_fd_sc_hd__inv_1 _08081_ (.A(_05617_),
    .Y(_02690_));
 sky130_fd_sc_hd__o311ai_4 _08082_ (.A1(_05621_),
    .A2(_02604_),
    .A3(_02605_),
    .B1(_02672_),
    .C1(_02666_),
    .Y(_02691_));
 sky130_fd_sc_hd__o21ai_2 _08083_ (.A1(_05660_),
    .A2(_02607_),
    .B1(_02529_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand4_1 _08084_ (.A(_02689_),
    .B(_02690_),
    .C(_02691_),
    .D(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__o211ai_1 _08085_ (.A1(_05687_),
    .A2(_02610_),
    .B1(_02523_),
    .C1(_02677_),
    .Y(_02694_));
 sky130_fd_sc_hd__a21oi_1 _08086_ (.A1(_02677_),
    .A2(_05696_),
    .B1(_05613_),
    .Y(_02695_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_02694_),
    .B(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__a31oi_1 _08088_ (.A1(_02687_),
    .A2(_02688_),
    .A3(_02693_),
    .B1(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__xnor2_1 _08089_ (.A(_05704_),
    .B(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__or3_1 _08090_ (.A(_05548_),
    .B(_05690_),
    .C(_05699_),
    .X(_02699_));
 sky130_fd_sc_hd__nor2_1 _08091_ (.A(_02628_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__a21boi_4 _08092_ (.A1(_02623_),
    .A2(_02627_),
    .B1_N(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__or2_0 _08093_ (.A(_05548_),
    .B(_05699_),
    .X(_02702_));
 sky130_fd_sc_hd__nor2_2 _08094_ (.A(_05548_),
    .B(_05699_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand3_1 _08095_ (.A(_02655_),
    .B(_02619_),
    .C(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nor2b_1 _08096_ (.A(_05548_),
    .B_N(_05700_),
    .Y(_02705_));
 sky130_fd_sc_hd__nor2_1 _08097_ (.A(_05549_),
    .B(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__o221ai_4 _08098_ (.A1(_02620_),
    .A2(_02702_),
    .B1(_02704_),
    .B2(_02618_),
    .C1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nor2_2 _08099_ (.A(_02701_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__xnor2_1 _08100_ (.A(_05708_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__o22ai_2 _08101_ (.A1(_02601_),
    .A2(_02698_),
    .B1(_02709_),
    .B2(_02632_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_1 _08102_ (.A(_01035_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__nor2_1 _08103_ (.A(\CPU_dmem_rd_data_a5[12] ),
    .B(_01036_),
    .Y(_02712_));
 sky130_fd_sc_hd__or3_4 _08104_ (.A(CPU_reset_a3),
    .B(_02711_),
    .C(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__nand3_1 _08110_ (.A(net1615),
    .B(net96),
    .C(_02596_),
    .Y(_02719_));
 sky130_fd_sc_hd__o21ai_0 _08111_ (.A1(_02596_),
    .A2(_02713_),
    .B1(_02719_),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_1 _08112_ (.A(_05704_),
    .Y(_02720_));
 sky130_fd_sc_hd__a21o_2 _08113_ (.A1(_05613_),
    .A2(_02720_),
    .B1(_05705_),
    .X(_02721_));
 sky130_fd_sc_hd__a21oi_1 _08114_ (.A1(_05617_),
    .A2(_02613_),
    .B1(_05678_),
    .Y(_02722_));
 sky130_fd_sc_hd__o21ai_1 _08115_ (.A1(_05669_),
    .A2(_02664_),
    .B1(_02603_),
    .Y(_02723_));
 sky130_fd_sc_hd__nor4_1 _08116_ (.A(_05612_),
    .B(_05686_),
    .C(_05695_),
    .D(_05704_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21boi_2 _08117_ (.A1(_02722_),
    .A2(_02723_),
    .B1_N(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _08118_ (.A(_02677_),
    .B(_02720_),
    .Y(_02726_));
 sky130_fd_sc_hd__nor2_1 _08119_ (.A(_02662_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__nor3_1 _08120_ (.A(_02721_),
    .B(_02725_),
    .C(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _08121_ (.A(_02603_),
    .B(_02724_),
    .Y(_02729_));
 sky130_fd_sc_hd__or2_0 _08122_ (.A(_02673_),
    .B(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__inv_1 _08123_ (.A(_05713_),
    .Y(_02731_));
 sky130_fd_sc_hd__a21oi_1 _08124_ (.A1(_02728_),
    .A2(_02730_),
    .B1(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__and3_1 _08125_ (.A(_02731_),
    .B(_02728_),
    .C(_02730_),
    .X(_02733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__o21ai_4 _08127_ (.A1(_02732_),
    .A2(_02733_),
    .B1(_02679_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor2_1 _08128_ (.A(_05708_),
    .B(_02699_),
    .Y(_02736_));
 sky130_fd_sc_hd__o21ai_1 _08129_ (.A1(_02652_),
    .A2(_02657_),
    .B1(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__nor2b_1 _08130_ (.A(_05699_),
    .B_N(_05691_),
    .Y(_02738_));
 sky130_fd_sc_hd__inv_1 _08131_ (.A(_05548_),
    .Y(_02739_));
 sky130_fd_sc_hd__o21a_1 _08132_ (.A1(_05700_),
    .A2(_02738_),
    .B1(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__inv_1 _08133_ (.A(_05708_),
    .Y(_02741_));
 sky130_fd_sc_hd__o21ai_0 _08134_ (.A1(_05549_),
    .A2(_02740_),
    .B1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__nor2b_1 _08135_ (.A(_05709_),
    .B_N(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__a21boi_1 _08136_ (.A1(_02737_),
    .A2(_02743_),
    .B1_N(_05717_),
    .Y(_02744_));
 sky130_fd_sc_hd__and3b_1 _08137_ (.A_N(_05717_),
    .B(_02737_),
    .C(_02743_),
    .X(_02745_));
 sky130_fd_sc_hd__o21ai_4 _08138_ (.A1(_02744_),
    .A2(_02745_),
    .B1(_02483_),
    .Y(_02746_));
 sky130_fd_sc_hd__nor2_1 _08139_ (.A(\CPU_dmem_rd_data_a5[13] ),
    .B(_01036_),
    .Y(_02747_));
 sky130_fd_sc_hd__a31oi_4 _08140_ (.A1(_01036_),
    .A2(_02735_),
    .A3(_02746_),
    .B1(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_1 _08141_ (.A(_02580_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _08142_ (.A(net1404),
    .B(_02596_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21oi_1 _08143_ (.A1(_02749_),
    .A2(_02750_),
    .B1(net109),
    .Y(_00548_));
 sky130_fd_sc_hd__nor2_1 _08144_ (.A(_05708_),
    .B(_05717_),
    .Y(_02751_));
 sky130_fd_sc_hd__nor2b_1 _08145_ (.A(_05717_),
    .B_N(_05709_),
    .Y(_02752_));
 sky130_fd_sc_hd__nor2_1 _08146_ (.A(_05718_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__o21ai_2 _08147_ (.A1(_05549_),
    .A2(_02705_),
    .B1(_02751_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_02753_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__a31oi_2 _08149_ (.A1(_02630_),
    .A2(_02703_),
    .A3(_02751_),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_2 _08150_ (.A(_01061_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__nor3_1 _08151_ (.A(_05668_),
    .B(_05713_),
    .C(_02729_),
    .Y(_02758_));
 sky130_fd_sc_hd__a2111oi_2 _08152_ (.A1(_02611_),
    .A2(_02614_),
    .B1(_02726_),
    .C1(_05713_),
    .D1(_05695_),
    .Y(_02759_));
 sky130_fd_sc_hd__a21oi_1 _08153_ (.A1(_05705_),
    .A2(_02731_),
    .B1(_05714_),
    .Y(_02760_));
 sky130_fd_sc_hd__o31ai_2 _08154_ (.A1(_05704_),
    .A2(_05713_),
    .A3(_02695_),
    .B1(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__a211oi_4 _08155_ (.A1(_02609_),
    .A2(_02758_),
    .B1(_02759_),
    .C1(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__xnor2_1 _08156_ (.A(_02543_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__a22oi_4 _08157_ (.A1(net98),
    .A2(_02757_),
    .B1(_02763_),
    .B2(_02679_),
    .Y(_02764_));
 sky130_fd_sc_hd__nor2_1 _08158_ (.A(\CPU_dmem_rd_data_a5[14] ),
    .B(_01036_),
    .Y(_02765_));
 sky130_fd_sc_hd__a211o_4 _08159_ (.A1(_01036_),
    .A2(_02764_),
    .B1(_02765_),
    .C1(net108),
    .X(_02766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_369 ();
 sky130_fd_sc_hd__nand3_1 _08161_ (.A(net1402),
    .B(net97),
    .C(_02596_),
    .Y(_02768_));
 sky130_fd_sc_hd__o21ai_0 _08162_ (.A1(_02596_),
    .A2(_02766_),
    .B1(_02768_),
    .Y(_00549_));
 sky130_fd_sc_hd__nor3_4 _08163_ (.A(_05708_),
    .B(_05717_),
    .C(_05726_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(_02739_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__a21oi_1 _08165_ (.A1(_05549_),
    .A2(_02741_),
    .B1(_05709_),
    .Y(_02771_));
 sky130_fd_sc_hd__a21oi_1 _08166_ (.A1(_05718_),
    .A2(_01061_),
    .B1(_05727_),
    .Y(_02772_));
 sky130_fd_sc_hd__o31ai_4 _08167_ (.A1(_05717_),
    .A2(_05726_),
    .A3(_02771_),
    .B1(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__inv_1 _08168_ (.A(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o31ai_1 _08169_ (.A1(_02646_),
    .A2(_02658_),
    .A3(_02770_),
    .B1(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__xor2_2 _08170_ (.A(_05543_),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__a21o_1 _08171_ (.A1(_05714_),
    .A2(_02543_),
    .B1(_05723_),
    .X(_02777_));
 sky130_fd_sc_hd__or2_1 _08172_ (.A(_05713_),
    .B(_05722_),
    .X(_02778_));
 sky130_fd_sc_hd__a21oi_1 _08173_ (.A1(_02728_),
    .A2(_02730_),
    .B1(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__or4_1 _08174_ (.A(_05608_),
    .B(_02601_),
    .C(_02777_),
    .D(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__o211ai_2 _08175_ (.A1(_02777_),
    .A2(_02779_),
    .B1(_05608_),
    .C1(_02679_),
    .Y(_02781_));
 sky130_fd_sc_hd__o211ai_4 _08176_ (.A1(_02632_),
    .A2(_02776_),
    .B1(_02780_),
    .C1(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2b_1 _08177_ (.A_N(\CPU_dmem_rd_data_a5[15] ),
    .B(_01035_),
    .Y(_02783_));
 sky130_fd_sc_hd__o211ai_4 _08178_ (.A1(_01035_),
    .A2(_02782_),
    .B1(_02783_),
    .C1(net97),
    .Y(_02784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_368 ();
 sky130_fd_sc_hd__nand3_1 _08180_ (.A(net1444),
    .B(net97),
    .C(_02596_),
    .Y(_02786_));
 sky130_fd_sc_hd__o21ai_0 _08181_ (.A1(_02596_),
    .A2(_02784_),
    .B1(_02786_),
    .Y(_00550_));
 sky130_fd_sc_hd__o21ai_0 _08182_ (.A1(_02701_),
    .A2(_02707_),
    .B1(_02769_),
    .Y(_02787_));
 sky130_fd_sc_hd__nor2b_1 _08183_ (.A(_05543_),
    .B_N(_05727_),
    .Y(_02788_));
 sky130_fd_sc_hd__nor2_1 _08184_ (.A(_05544_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__nor2_1 _08185_ (.A(_05543_),
    .B(_05726_),
    .Y(_02790_));
 sky130_fd_sc_hd__o21ai_0 _08186_ (.A1(_05718_),
    .A2(_02752_),
    .B1(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__and2_0 _08187_ (.A(_02789_),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__o21ai_1 _08188_ (.A1(_05543_),
    .A2(_02787_),
    .B1(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__inv_1 _08189_ (.A(_05730_),
    .Y(_02794_));
 sky130_fd_sc_hd__nor2_1 _08190_ (.A(_02794_),
    .B(_02632_),
    .Y(_02795_));
 sky130_fd_sc_hd__inv_1 _08191_ (.A(_05604_),
    .Y(_02796_));
 sky130_fd_sc_hd__inv_1 _08192_ (.A(_05608_),
    .Y(_02797_));
 sky130_fd_sc_hd__a21oi_1 _08193_ (.A1(_02797_),
    .A2(_05723_),
    .B1(_05609_),
    .Y(_02798_));
 sky130_fd_sc_hd__o31ai_1 _08194_ (.A1(_05608_),
    .A2(_05722_),
    .A3(_02760_),
    .B1(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__nor4_1 _08195_ (.A(_05608_),
    .B(_05704_),
    .C(_05713_),
    .D(_05722_),
    .Y(_02800_));
 sky130_fd_sc_hd__nand3_1 _08196_ (.A(_02687_),
    .B(_02688_),
    .C(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__a41oi_4 _08197_ (.A1(_02689_),
    .A2(_02690_),
    .A3(_02691_),
    .A4(_02692_),
    .B1(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__a21boi_1 _08198_ (.A1(_02694_),
    .A2(_02695_),
    .B1_N(_02800_),
    .Y(_02803_));
 sky130_fd_sc_hd__nor3_1 _08199_ (.A(_02799_),
    .B(_02802_),
    .C(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__xnor2_1 _08200_ (.A(_02796_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o2111a_1 _08201_ (.A1(_05543_),
    .A2(_02787_),
    .B1(_02792_),
    .C1(net98),
    .D1(_02794_),
    .X(_02806_));
 sky130_fd_sc_hd__a221oi_4 _08202_ (.A1(_02793_),
    .A2(_02795_),
    .B1(_02805_),
    .B2(_02679_),
    .C1(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _08203_ (.A(_01036_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__o211ai_4 _08204_ (.A1(\CPU_dmem_rd_data_a5[16] ),
    .A2(_01036_),
    .B1(_02808_),
    .C1(net97),
    .Y(_02809_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_367 ();
 sky130_fd_sc_hd__nand3_1 _08206_ (.A(net1447),
    .B(net97),
    .C(_02596_),
    .Y(_02811_));
 sky130_fd_sc_hd__o21ai_0 _08207_ (.A1(_02596_),
    .A2(_02809_),
    .B1(_02811_),
    .Y(_00551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_366 ();
 sky130_fd_sc_hd__a21oi_1 _08209_ (.A1(_05544_),
    .A2(_02794_),
    .B1(_05731_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21bo_1 _08210_ (.A1(_02740_),
    .A2(_02769_),
    .B1_N(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__nor2_1 _08211_ (.A(_02773_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__nor2b_1 _08212_ (.A(_02699_),
    .B_N(_02769_),
    .Y(_02816_));
 sky130_fd_sc_hd__and3_1 _08213_ (.A(_02624_),
    .B(_02700_),
    .C(_02769_),
    .X(_02817_));
 sky130_fd_sc_hd__nand2_2 _08214_ (.A(_02649_),
    .B(_02651_),
    .Y(_02818_));
 sky130_fd_sc_hd__a22oi_4 _08215_ (.A1(_02657_),
    .A2(_02816_),
    .B1(_02817_),
    .B2(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2b_1 _08216_ (.A_N(_05544_),
    .B(_05543_),
    .Y(_02820_));
 sky130_fd_sc_hd__a21oi_1 _08217_ (.A1(_02794_),
    .A2(_02820_),
    .B1(_05731_),
    .Y(_02821_));
 sky130_fd_sc_hd__a21oi_1 _08218_ (.A1(_02815_),
    .A2(_02819_),
    .B1(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__xnor2_2 _08219_ (.A(_05734_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__inv_1 _08220_ (.A(_05599_),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _08221_ (.A(_02728_),
    .B(_02730_),
    .Y(_02825_));
 sky130_fd_sc_hd__nor3_2 _08222_ (.A(_05604_),
    .B(_05608_),
    .C(_02778_),
    .Y(_02826_));
 sky130_fd_sc_hd__a21oi_2 _08223_ (.A1(_05714_),
    .A2(_02543_),
    .B1(_05723_),
    .Y(_02827_));
 sky130_fd_sc_hd__a21oi_2 _08224_ (.A1(_02796_),
    .A2(_05609_),
    .B1(_05605_),
    .Y(_02828_));
 sky130_fd_sc_hd__o31ai_2 _08225_ (.A1(_05604_),
    .A2(_05608_),
    .A3(_02827_),
    .B1(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__a21oi_1 _08226_ (.A1(_02825_),
    .A2(_02826_),
    .B1(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__xnor2_1 _08227_ (.A(_02824_),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__a22oi_4 _08228_ (.A1(net98),
    .A2(_02823_),
    .B1(_02831_),
    .B2(_02679_),
    .Y(_02832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_365 ();
 sky130_fd_sc_hd__nand3_4 _08230_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[17] ),
    .C(_01035_),
    .Y(_02834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_363 ();
 sky130_fd_sc_hd__nand3_1 _08233_ (.A(net1573),
    .B(net97),
    .C(_02596_),
    .Y(_02837_));
 sky130_fd_sc_hd__o221ai_1 _08234_ (.A1(_02582_),
    .A2(_02832_),
    .B1(_02834_),
    .B2(_02596_),
    .C1(_02837_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand4_1 _08235_ (.A(_02824_),
    .B(_02796_),
    .C(_02797_),
    .D(_02543_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21oi_1 _08236_ (.A1(_02824_),
    .A2(_05605_),
    .B1(_05600_),
    .Y(_02839_));
 sky130_fd_sc_hd__o31ai_1 _08237_ (.A1(_05599_),
    .A2(_05604_),
    .A3(_02798_),
    .B1(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__o21bai_1 _08238_ (.A1(_02762_),
    .A2(_02838_),
    .B1_N(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__xnor2_1 _08239_ (.A(_05739_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__inv_1 _08240_ (.A(_05743_),
    .Y(_02843_));
 sky130_fd_sc_hd__nor2_1 _08241_ (.A(_05730_),
    .B(_05734_),
    .Y(_02844_));
 sky130_fd_sc_hd__and4_1 _08242_ (.A(_02703_),
    .B(_02751_),
    .C(_02790_),
    .D(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__o31ai_2 _08243_ (.A1(_05544_),
    .A2(_02788_),
    .A3(_02790_),
    .B1(_02844_),
    .Y(_02846_));
 sky130_fd_sc_hd__a31oi_4 _08244_ (.A1(_02753_),
    .A2(_02754_),
    .A3(_02789_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__inv_1 _08245_ (.A(_05734_),
    .Y(_02848_));
 sky130_fd_sc_hd__a21oi_2 _08246_ (.A1(_05731_),
    .A2(_02848_),
    .B1(_05735_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2b_1 _08247_ (.A_N(_02847_),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__a21oi_1 _08248_ (.A1(_02630_),
    .A2(_02845_),
    .B1(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__xnor2_2 _08249_ (.A(_02843_),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__a22oi_4 _08250_ (.A1(_02679_),
    .A2(_02842_),
    .B1(_02852_),
    .B2(net98),
    .Y(_02853_));
 sky130_fd_sc_hd__nand2_4 _08251_ (.A(_01036_),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__nor2_4 _08252_ (.A(\CPU_dmem_rd_data_a5[18] ),
    .B(_01036_),
    .Y(_02855_));
 sky130_fd_sc_hd__nor2_8 _08253_ (.A(net108),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_362 ();
 sky130_fd_sc_hd__and3_1 _08255_ (.A(net1835),
    .B(_02586_),
    .C(_02596_),
    .X(_02858_));
 sky130_fd_sc_hd__a31o_1 _08256_ (.A1(_02580_),
    .A2(_02854_),
    .A3(_02856_),
    .B1(_02858_),
    .X(_00553_));
 sky130_fd_sc_hd__or4_1 _08257_ (.A(_05543_),
    .B(_05730_),
    .C(_05734_),
    .D(_05743_),
    .X(_02859_));
 sky130_fd_sc_hd__nor4_1 _08258_ (.A(_05543_),
    .B(_05730_),
    .C(_05734_),
    .D(_05743_),
    .Y(_02860_));
 sky130_fd_sc_hd__a21oi_1 _08259_ (.A1(_05735_),
    .A2(_02843_),
    .B1(_05744_),
    .Y(_02861_));
 sky130_fd_sc_hd__o31ai_1 _08260_ (.A1(_05734_),
    .A2(_05743_),
    .A3(_02813_),
    .B1(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__a21oi_1 _08261_ (.A1(_02773_),
    .A2(_02860_),
    .B1(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__o41ai_1 _08262_ (.A1(_02646_),
    .A2(_02658_),
    .A3(_02770_),
    .A4(_02859_),
    .B1(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__xnor2_1 _08263_ (.A(_01065_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__nor2_4 _08264_ (.A(_02632_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__inv_1 _08265_ (.A(_05594_),
    .Y(_02867_));
 sky130_fd_sc_hd__a211o_1 _08266_ (.A1(_02665_),
    .A2(_02673_),
    .B1(_02729_),
    .C1(_02778_),
    .X(_02868_));
 sky130_fd_sc_hd__nor2_1 _08267_ (.A(_05713_),
    .B(_05722_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_1 _08268_ (.A(_02726_),
    .B(_02778_),
    .Y(_02870_));
 sky130_fd_sc_hd__o21ai_2 _08269_ (.A1(_02722_),
    .A2(_02675_),
    .B1(_02662_),
    .Y(_02871_));
 sky130_fd_sc_hd__a21oi_4 _08270_ (.A1(_05600_),
    .A2(_02499_),
    .B1(_05740_),
    .Y(_02872_));
 sky130_fd_sc_hd__o311ai_4 _08271_ (.A1(_05599_),
    .A2(_05739_),
    .A3(_02828_),
    .B1(_02872_),
    .C1(_02827_),
    .Y(_02873_));
 sky130_fd_sc_hd__a221oi_4 _08272_ (.A1(_02721_),
    .A2(_02869_),
    .B1(_02870_),
    .B2(_02871_),
    .C1(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand2b_1 _08273_ (.A_N(_05609_),
    .B(_05608_),
    .Y(_02875_));
 sky130_fd_sc_hd__a21oi_1 _08274_ (.A1(_02796_),
    .A2(_02875_),
    .B1(_05605_),
    .Y(_02876_));
 sky130_fd_sc_hd__o21bai_1 _08275_ (.A1(_05599_),
    .A2(_02876_),
    .B1_N(_05600_),
    .Y(_02877_));
 sky130_fd_sc_hd__a21oi_1 _08276_ (.A1(_02499_),
    .A2(_02877_),
    .B1(_05740_),
    .Y(_02878_));
 sky130_fd_sc_hd__a21oi_1 _08277_ (.A1(_02868_),
    .A2(_02874_),
    .B1(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__xnor2_1 _08278_ (.A(_02867_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__nor2_2 _08279_ (.A(_02601_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__nor2_8 _08280_ (.A(_02866_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_361 ();
 sky130_fd_sc_hd__and3_4 _08282_ (.A(_02586_),
    .B(\CPU_dmem_rd_data_a5[19] ),
    .C(_01035_),
    .X(_02884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_360 ();
 sky130_fd_sc_hd__and3_1 _08284_ (.A(net1751),
    .B(net97),
    .C(_02596_),
    .X(_02886_));
 sky130_fd_sc_hd__a21oi_1 _08285_ (.A1(_02580_),
    .A2(_02884_),
    .B1(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21ai_0 _08286_ (.A1(_02582_),
    .A2(_02882_),
    .B1(_02887_),
    .Y(_00554_));
 sky130_fd_sc_hd__a22o_2 _08287_ (.A1(_05518_),
    .A2(_02483_),
    .B1(_02679_),
    .B2(_05514_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2i_4 _08288_ (.A0(\CPU_dmem_rd_data_a5[1] ),
    .A1(_02888_),
    .S(_01036_),
    .Y(_02889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_359 ();
 sky130_fd_sc_hd__nand2_1 _08290_ (.A(net1434),
    .B(_02596_),
    .Y(_02891_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_357 ();
 sky130_fd_sc_hd__o211ai_1 _08293_ (.A1(_02596_),
    .A2(_02889_),
    .B1(_02891_),
    .C1(_02586_),
    .Y(_00555_));
 sky130_fd_sc_hd__nor4_1 _08294_ (.A(_05594_),
    .B(_05599_),
    .C(_05604_),
    .D(_05739_),
    .Y(_02894_));
 sky130_fd_sc_hd__o31ai_2 _08295_ (.A1(_02799_),
    .A2(_02802_),
    .A3(_02803_),
    .B1(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__o21bai_1 _08296_ (.A1(_05739_),
    .A2(_02839_),
    .B1_N(_05740_),
    .Y(_02896_));
 sky130_fd_sc_hd__a21oi_1 _08297_ (.A1(_02867_),
    .A2(_02896_),
    .B1(_05595_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_2 _08298_ (.A(_02895_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__xnor2_1 _08299_ (.A(_05748_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _08300_ (.A(_02769_),
    .B(_02860_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand3_1 _08301_ (.A(_01065_),
    .B(_02843_),
    .C(_02844_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21oi_1 _08302_ (.A1(_02789_),
    .A2(_02791_),
    .B1(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a21oi_1 _08303_ (.A1(_01065_),
    .A2(_05744_),
    .B1(_05539_),
    .Y(_02903_));
 sky130_fd_sc_hd__o31ai_1 _08304_ (.A1(_05538_),
    .A2(_05743_),
    .A3(_02849_),
    .B1(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nor2_1 _08305_ (.A(_02902_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__o31ai_4 _08306_ (.A1(_05538_),
    .A2(_02708_),
    .A3(_02900_),
    .B1(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__xnor2_2 _08307_ (.A(_05752_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__a22oi_4 _08308_ (.A1(_02679_),
    .A2(_02899_),
    .B1(_02907_),
    .B2(net98),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_4 _08309_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[20] ),
    .C(_01035_),
    .Y(_02909_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_356 ();
 sky130_fd_sc_hd__nand3_1 _08311_ (.A(net1505),
    .B(net96),
    .C(_02596_),
    .Y(_02911_));
 sky130_fd_sc_hd__o221ai_1 _08312_ (.A1(_02582_),
    .A2(_02908_),
    .B1(_02909_),
    .B2(_02596_),
    .C1(_02911_),
    .Y(_00556_));
 sky130_fd_sc_hd__a21oi_1 _08313_ (.A1(_05539_),
    .A2(_01066_),
    .B1(_05753_),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _08314_ (.A(_02861_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__nor3_2 _08315_ (.A(_02773_),
    .B(_02814_),
    .C(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__o31a_1 _08316_ (.A1(_05734_),
    .A2(_05743_),
    .A3(_02821_),
    .B1(_02861_),
    .X(_02915_));
 sky130_fd_sc_hd__o31a_1 _08317_ (.A1(_05538_),
    .A2(_05752_),
    .A3(_02915_),
    .B1(_02912_),
    .X(_02916_));
 sky130_fd_sc_hd__a211oi_4 _08318_ (.A1(_02819_),
    .A2(_02914_),
    .B1(_02916_),
    .C1(_05761_),
    .Y(_02917_));
 sky130_fd_sc_hd__inv_1 _08319_ (.A(_05761_),
    .Y(_02918_));
 sky130_fd_sc_hd__a21oi_1 _08320_ (.A1(_02819_),
    .A2(_02914_),
    .B1(_02916_),
    .Y(_02919_));
 sky130_fd_sc_hd__nor2_1 _08321_ (.A(_02918_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__nor2b_1 _08322_ (.A(_05748_),
    .B_N(_05595_),
    .Y(_02921_));
 sky130_fd_sc_hd__nor2_1 _08323_ (.A(_05749_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__o31ai_4 _08324_ (.A1(_05594_),
    .A2(_05748_),
    .A3(_02872_),
    .B1(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__nor2_1 _08325_ (.A(_05594_),
    .B(_05748_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2b_1 _08326_ (.A_N(_05740_),
    .B(_05739_),
    .Y(_02925_));
 sky130_fd_sc_hd__or3b_1 _08327_ (.A(_05600_),
    .B(_05740_),
    .C_N(_05599_),
    .X(_02926_));
 sky130_fd_sc_hd__a311o_2 _08328_ (.A1(_02924_),
    .A2(_02925_),
    .A3(_02926_),
    .B1(_02921_),
    .C1(_05749_),
    .X(_02927_));
 sky130_fd_sc_hd__o311ai_4 _08329_ (.A1(_02721_),
    .A2(_02725_),
    .A3(_02727_),
    .B1(_02826_),
    .C1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand4_1 _08330_ (.A(_02603_),
    .B(_02724_),
    .C(_02826_),
    .D(_02927_),
    .Y(_02929_));
 sky130_fd_sc_hd__a2bb2oi_2 _08331_ (.A1_N(_02673_),
    .A2_N(_02929_),
    .B1(_02927_),
    .B2(_02829_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand2_1 _08332_ (.A(_02928_),
    .B(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__nor2_1 _08333_ (.A(_02923_),
    .B(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__xnor2_1 _08334_ (.A(_05757_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__o32a_4 _08335_ (.A1(_02632_),
    .A2(_02917_),
    .A3(_02920_),
    .B1(_02601_),
    .B2(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_355 ();
 sky130_fd_sc_hd__nand3_4 _08337_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[21] ),
    .C(_01035_),
    .Y(_02936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_354 ();
 sky130_fd_sc_hd__nand3_1 _08339_ (.A(net1649),
    .B(_02586_),
    .C(_02596_),
    .Y(_02938_));
 sky130_fd_sc_hd__o221ai_1 _08340_ (.A1(_02582_),
    .A2(_02934_),
    .B1(_02936_),
    .B2(_02596_),
    .C1(_02938_),
    .Y(_00557_));
 sky130_fd_sc_hd__nor4_1 _08341_ (.A(_05594_),
    .B(_05739_),
    .C(_05748_),
    .D(_05757_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2b_1 _08342_ (.A_N(_02838_),
    .B(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__a21oi_1 _08343_ (.A1(_02867_),
    .A2(_05740_),
    .B1(_05595_),
    .Y(_02941_));
 sky130_fd_sc_hd__nor2b_1 _08344_ (.A(_05757_),
    .B_N(_05749_),
    .Y(_02942_));
 sky130_fd_sc_hd__nor2_1 _08345_ (.A(_05758_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__o31ai_1 _08346_ (.A1(_05748_),
    .A2(_05757_),
    .A3(_02941_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__a21oi_1 _08347_ (.A1(_02840_),
    .A2(_02939_),
    .B1(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__o21ai_4 _08348_ (.A1(_02762_),
    .A2(_02940_),
    .B1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__xnor2_1 _08349_ (.A(_05766_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__or2_2 _08350_ (.A(_05752_),
    .B(_05761_),
    .X(_02948_));
 sky130_fd_sc_hd__a21oi_2 _08351_ (.A1(_05753_),
    .A2(_02918_),
    .B1(_05762_),
    .Y(_02949_));
 sky130_fd_sc_hd__o211ai_1 _08352_ (.A1(_02903_),
    .A2(_02948_),
    .B1(_02949_),
    .C1(_02849_),
    .Y(_02950_));
 sky130_fd_sc_hd__nor4_2 _08353_ (.A(_02621_),
    .B(_02629_),
    .C(_02847_),
    .D(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__nand4_1 _08354_ (.A(_02703_),
    .B(_02751_),
    .C(_02790_),
    .D(_02844_),
    .Y(_02952_));
 sky130_fd_sc_hd__o2111ai_1 _08355_ (.A1(_02903_),
    .A2(_02948_),
    .B1(_02949_),
    .C1(_02849_),
    .D1(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__or3_1 _08356_ (.A(_05538_),
    .B(_05743_),
    .C(_02948_),
    .X(_02954_));
 sky130_fd_sc_hd__o211ai_1 _08357_ (.A1(_02903_),
    .A2(_02948_),
    .B1(_02954_),
    .C1(_02949_),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ai_2 _08358_ (.A1(_02847_),
    .A2(_02953_),
    .B1(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__nor2_1 _08359_ (.A(_02951_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__xnor2_2 _08360_ (.A(_05770_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__a22oi_4 _08361_ (.A1(_02679_),
    .A2(_02947_),
    .B1(_02958_),
    .B2(_02483_),
    .Y(_02959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_353 ();
 sky130_fd_sc_hd__and3_4 _08363_ (.A(_02586_),
    .B(\CPU_dmem_rd_data_a5[22] ),
    .C(_01035_),
    .X(_02961_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_352 ();
 sky130_fd_sc_hd__and3_1 _08365_ (.A(net1818),
    .B(_02586_),
    .C(_02596_),
    .X(_02963_));
 sky130_fd_sc_hd__a21oi_1 _08366_ (.A1(_02580_),
    .A2(_02961_),
    .B1(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__o21ai_0 _08367_ (.A1(_02582_),
    .A2(_02959_),
    .B1(_02964_),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_1 _08368_ (.A(_05590_),
    .Y(_02965_));
 sky130_fd_sc_hd__inv_1 _08369_ (.A(_05757_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_2 _08370_ (.A(_02966_),
    .B(_02512_),
    .Y(_02967_));
 sky130_fd_sc_hd__a21oi_1 _08371_ (.A1(_05758_),
    .A2(_02512_),
    .B1(_05767_),
    .Y(_02968_));
 sky130_fd_sc_hd__o21ai_0 _08372_ (.A1(_02922_),
    .A2(_02967_),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand3_1 _08373_ (.A(_02966_),
    .B(_02512_),
    .C(_02924_),
    .Y(_02970_));
 sky130_fd_sc_hd__a211oi_2 _08374_ (.A1(_02868_),
    .A2(_02874_),
    .B1(_02970_),
    .C1(_02878_),
    .Y(_02971_));
 sky130_fd_sc_hd__nor2_1 _08375_ (.A(_02969_),
    .B(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__xnor2_1 _08376_ (.A(_02965_),
    .B(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__or3_1 _08377_ (.A(_05538_),
    .B(_05770_),
    .C(_02948_),
    .X(_02974_));
 sky130_fd_sc_hd__inv_1 _08378_ (.A(_05770_),
    .Y(_02975_));
 sky130_fd_sc_hd__a21oi_1 _08379_ (.A1(_05762_),
    .A2(_02975_),
    .B1(_05771_),
    .Y(_02976_));
 sky130_fd_sc_hd__o31a_1 _08380_ (.A1(_05761_),
    .A2(_05770_),
    .A3(_02912_),
    .B1(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__o21a_1 _08381_ (.A1(_02863_),
    .A2(_02974_),
    .B1(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__or2_0 _08382_ (.A(_02900_),
    .B(_02974_),
    .X(_02979_));
 sky130_fd_sc_hd__or4_2 _08383_ (.A(_05548_),
    .B(_02646_),
    .C(_02658_),
    .D(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(_02978_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__xnor2_2 _08385_ (.A(_05533_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__a22oi_4 _08386_ (.A1(_02679_),
    .A2(_02973_),
    .B1(_02982_),
    .B2(net98),
    .Y(_02983_));
 sky130_fd_sc_hd__nand3_4 _08387_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[23] ),
    .C(_01035_),
    .Y(_02984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_351 ();
 sky130_fd_sc_hd__nand3_1 _08389_ (.A(net1519),
    .B(_02586_),
    .C(_02596_),
    .Y(_02986_));
 sky130_fd_sc_hd__o221ai_1 _08390_ (.A1(_02582_),
    .A2(_02983_),
    .B1(_02984_),
    .B2(_02596_),
    .C1(_02986_),
    .Y(_00559_));
 sky130_fd_sc_hd__inv_1 _08391_ (.A(_05586_),
    .Y(_02987_));
 sky130_fd_sc_hd__nor2_1 _08392_ (.A(_02987_),
    .B(_02601_),
    .Y(_02988_));
 sky130_fd_sc_hd__nor2_1 _08393_ (.A(_05586_),
    .B(_02601_),
    .Y(_02989_));
 sky130_fd_sc_hd__inv_1 _08394_ (.A(_05767_),
    .Y(_02990_));
 sky130_fd_sc_hd__o21ai_0 _08395_ (.A1(_05758_),
    .A2(_02942_),
    .B1(_02512_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21oi_1 _08396_ (.A1(_02990_),
    .A2(_02991_),
    .B1(_05590_),
    .Y(_02992_));
 sky130_fd_sc_hd__nor2_2 _08397_ (.A(_05591_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__nor3_1 _08398_ (.A(_05590_),
    .B(_05748_),
    .C(_02967_),
    .Y(_02994_));
 sky130_fd_sc_hd__nor3_1 _08399_ (.A(_05591_),
    .B(_02992_),
    .C(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__a31o_1 _08400_ (.A1(_02895_),
    .A2(_02897_),
    .A3(_02993_),
    .B1(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2i_4 _08401_ (.A0(_02988_),
    .A1(_02989_),
    .S(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__o21ba_1 _08402_ (.A1(_05770_),
    .A2(_02949_),
    .B1_N(_05771_),
    .X(_02998_));
 sky130_fd_sc_hd__o21ba_1 _08403_ (.A1(_05533_),
    .A2(_02998_),
    .B1_N(_05534_),
    .X(_02999_));
 sky130_fd_sc_hd__nor3_2 _08404_ (.A(_05533_),
    .B(_05770_),
    .C(_02948_),
    .Y(_03000_));
 sky130_fd_sc_hd__and3_1 _08405_ (.A(_01065_),
    .B(_02860_),
    .C(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__o211ai_2 _08406_ (.A1(_02701_),
    .A2(_02707_),
    .B1(_02769_),
    .C1(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__o21ai_1 _08407_ (.A1(_02902_),
    .A2(_02904_),
    .B1(_03000_),
    .Y(_03003_));
 sky130_fd_sc_hd__inv_1 _08408_ (.A(_05774_),
    .Y(_03004_));
 sky130_fd_sc_hd__a31o_1 _08409_ (.A1(_02999_),
    .A2(_03002_),
    .A3(_03003_),
    .B1(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__nand4_1 _08410_ (.A(_03004_),
    .B(_02999_),
    .C(_03002_),
    .D(_03003_),
    .Y(_03006_));
 sky130_fd_sc_hd__a21o_2 _08411_ (.A1(_03005_),
    .A2(_03006_),
    .B1(_02632_),
    .X(_03007_));
 sky130_fd_sc_hd__nor2_1 _08412_ (.A(\CPU_dmem_rd_data_a5[24] ),
    .B(_01036_),
    .Y(_03008_));
 sky130_fd_sc_hd__a31oi_4 _08413_ (.A1(_01036_),
    .A2(_02997_),
    .A3(_03007_),
    .B1(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_1 _08414_ (.A(_02580_),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _08415_ (.A(net1405),
    .B(_02596_),
    .Y(_03011_));
 sky130_fd_sc_hd__a21oi_1 _08416_ (.A1(_03010_),
    .A2(_03011_),
    .B1(net109),
    .Y(_00560_));
 sky130_fd_sc_hd__o21bai_1 _08417_ (.A1(_05590_),
    .A2(_02968_),
    .B1_N(_05591_),
    .Y(_03012_));
 sky130_fd_sc_hd__a21oi_2 _08418_ (.A1(_02987_),
    .A2(_03012_),
    .B1(_05587_),
    .Y(_03013_));
 sky130_fd_sc_hd__o31ai_1 _08419_ (.A1(_05586_),
    .A2(_05590_),
    .A3(_02967_),
    .B1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand4b_1 _08420_ (.A_N(_02923_),
    .B(_02928_),
    .C(_02930_),
    .D(_03013_),
    .Y(_03015_));
 sky130_fd_sc_hd__and3_1 _08421_ (.A(_05581_),
    .B(_03014_),
    .C(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__a21oi_1 _08422_ (.A1(_03014_),
    .A2(_03015_),
    .B1(_05581_),
    .Y(_03017_));
 sky130_fd_sc_hd__o21ai_4 _08423_ (.A1(_03016_),
    .A2(_03017_),
    .B1(_02679_),
    .Y(_03018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_350 ();
 sky130_fd_sc_hd__inv_1 _08425_ (.A(_05778_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _08426_ (.A(_03020_),
    .B(_02632_),
    .Y(_03021_));
 sky130_fd_sc_hd__nor2_1 _08427_ (.A(_05778_),
    .B(_02632_),
    .Y(_03022_));
 sky130_fd_sc_hd__o21bai_1 _08428_ (.A1(_05533_),
    .A2(_02976_),
    .B1_N(_05534_),
    .Y(_03023_));
 sky130_fd_sc_hd__nor3_2 _08429_ (.A(_05533_),
    .B(_05770_),
    .C(_05774_),
    .Y(_03024_));
 sky130_fd_sc_hd__a221oi_4 _08430_ (.A1(_03004_),
    .A2(_03023_),
    .B1(_03024_),
    .B2(_02917_),
    .C1(_05775_),
    .Y(_03025_));
 sky130_fd_sc_hd__mux2i_4 _08431_ (.A0(_03021_),
    .A1(_03022_),
    .S(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_347 ();
 sky130_fd_sc_hd__nor2_1 _08435_ (.A(_01035_),
    .B(_02596_),
    .Y(_03030_));
 sky130_fd_sc_hd__nor2_8 _08436_ (.A(\CPU_dmem_rd_data_a5[25] ),
    .B(_01036_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(_02580_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__o21ai_0 _08438_ (.A1(net1722),
    .A2(_02580_),
    .B1(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_346 ();
 sky130_fd_sc_hd__a311oi_1 _08440_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03030_),
    .B1(_03033_),
    .C1(net108),
    .Y(_00561_));
 sky130_fd_sc_hd__nor2_1 _08441_ (.A(_05787_),
    .B(_02632_),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2_1 _08442_ (.A(_01046_),
    .B(_02632_),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _08443_ (.A(_03020_),
    .B(_03024_),
    .Y(_03037_));
 sky130_fd_sc_hd__a21oi_1 _08444_ (.A1(_01097_),
    .A2(_05771_),
    .B1(_05534_),
    .Y(_03038_));
 sky130_fd_sc_hd__o21bai_1 _08445_ (.A1(_05774_),
    .A2(_03038_),
    .B1_N(_05775_),
    .Y(_03039_));
 sky130_fd_sc_hd__a21oi_1 _08446_ (.A1(_03020_),
    .A2(_03039_),
    .B1(_05779_),
    .Y(_03040_));
 sky130_fd_sc_hd__o31ai_2 _08447_ (.A1(_02951_),
    .A2(_02956_),
    .A3(_03037_),
    .B1(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__mux2i_4 _08448_ (.A0(_03035_),
    .A1(_03036_),
    .S(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__inv_1 _08449_ (.A(_05581_),
    .Y(_03043_));
 sky130_fd_sc_hd__a21oi_1 _08450_ (.A1(_02965_),
    .A2(_05767_),
    .B1(_05591_),
    .Y(_03044_));
 sky130_fd_sc_hd__inv_1 _08451_ (.A(_05587_),
    .Y(_03045_));
 sky130_fd_sc_hd__o21ai_1 _08452_ (.A1(_05586_),
    .A2(_03044_),
    .B1(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__a21o_1 _08453_ (.A1(_03043_),
    .A2(_03046_),
    .B1(_05582_),
    .X(_03047_));
 sky130_fd_sc_hd__nor4_1 _08454_ (.A(_05581_),
    .B(_05586_),
    .C(_05590_),
    .D(_05766_),
    .Y(_03048_));
 sky130_fd_sc_hd__or2_0 _08455_ (.A(_03047_),
    .B(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__o2111ai_4 _08456_ (.A1(_02946_),
    .A2(_03047_),
    .B1(_03049_),
    .C1(_02679_),
    .D1(_05783_),
    .Y(_03050_));
 sky130_fd_sc_hd__a2111o_1 _08457_ (.A1(_02946_),
    .A2(_03048_),
    .B1(_03047_),
    .C1(_05783_),
    .D1(_02601_),
    .X(_03051_));
 sky130_fd_sc_hd__nor2_1 _08458_ (.A(\CPU_dmem_rd_data_a5[26] ),
    .B(_01036_),
    .Y(_03052_));
 sky130_fd_sc_hd__a41oi_4 _08459_ (.A1(_01036_),
    .A2(_03042_),
    .A3(_03050_),
    .A4(_03051_),
    .B1(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_1 _08460_ (.A(_02580_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _08461_ (.A(net1473),
    .B(_02596_),
    .Y(_03055_));
 sky130_fd_sc_hd__a21oi_1 _08462_ (.A1(_03054_),
    .A2(_03055_),
    .B1(net109),
    .Y(_00562_));
 sky130_fd_sc_hd__nor4_2 _08463_ (.A(_05581_),
    .B(_05586_),
    .C(_05590_),
    .D(_05783_),
    .Y(_03056_));
 sky130_fd_sc_hd__a2111oi_0 _08464_ (.A1(_02965_),
    .A2(_02969_),
    .B1(_05582_),
    .C1(_05587_),
    .D1(_05591_),
    .Y(_03057_));
 sky130_fd_sc_hd__a21oi_1 _08465_ (.A1(_05586_),
    .A2(_03045_),
    .B1(_05581_),
    .Y(_03058_));
 sky130_fd_sc_hd__nor2_1 _08466_ (.A(_05582_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__inv_1 _08467_ (.A(_05784_),
    .Y(_03060_));
 sky130_fd_sc_hd__o31a_1 _08468_ (.A1(_05783_),
    .A2(_03057_),
    .A3(_03059_),
    .B1(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__a21boi_0 _08469_ (.A1(_02971_),
    .A2(_03056_),
    .B1_N(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_1 _08470_ (.A(_05576_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21oi_1 _08471_ (.A1(_05534_),
    .A2(_03004_),
    .B1(_05775_),
    .Y(_03064_));
 sky130_fd_sc_hd__a21oi_2 _08472_ (.A1(_05779_),
    .A2(_01046_),
    .B1(_05788_),
    .Y(_03065_));
 sky130_fd_sc_hd__o31ai_2 _08473_ (.A1(_05778_),
    .A2(_05787_),
    .A3(_03064_),
    .B1(_03065_),
    .Y(_03066_));
 sky130_fd_sc_hd__nor4_2 _08474_ (.A(_05533_),
    .B(_05774_),
    .C(_05778_),
    .D(_05787_),
    .Y(_03067_));
 sky130_fd_sc_hd__nor4_1 _08475_ (.A(_05528_),
    .B(_02632_),
    .C(_03066_),
    .D(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__a31oi_1 _08476_ (.A1(_05528_),
    .A2(_02483_),
    .A3(_03066_),
    .B1(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__nor3_1 _08477_ (.A(_05528_),
    .B(_02632_),
    .C(_03066_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand3_1 _08478_ (.A(_05528_),
    .B(_02483_),
    .C(_03067_),
    .Y(_03071_));
 sky130_fd_sc_hd__a21oi_1 _08479_ (.A1(_02978_),
    .A2(_02980_),
    .B1(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__a31oi_1 _08480_ (.A1(_02978_),
    .A2(_02980_),
    .A3(_03070_),
    .B1(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__o211a_4 _08481_ (.A1(_02601_),
    .A2(_03063_),
    .B1(_03069_),
    .C1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_345 ();
 sky130_fd_sc_hd__nand3_4 _08483_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[27] ),
    .C(_01035_),
    .Y(_03076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_344 ();
 sky130_fd_sc_hd__nand3_1 _08485_ (.A(net1515),
    .B(net97),
    .C(_02596_),
    .Y(_03078_));
 sky130_fd_sc_hd__o221ai_1 _08486_ (.A1(_02582_),
    .A2(_03074_),
    .B1(_03076_),
    .B2(_02596_),
    .C1(_03078_),
    .Y(_00563_));
 sky130_fd_sc_hd__or4_2 _08487_ (.A(_05576_),
    .B(_05581_),
    .C(_05586_),
    .D(_05783_),
    .X(_03079_));
 sky130_fd_sc_hd__a21o_1 _08488_ (.A1(_03043_),
    .A2(_05587_),
    .B1(_05582_),
    .X(_03080_));
 sky130_fd_sc_hd__a21oi_2 _08489_ (.A1(_02516_),
    .A2(_03080_),
    .B1(_05784_),
    .Y(_03081_));
 sky130_fd_sc_hd__inv_1 _08490_ (.A(_05577_),
    .Y(_03082_));
 sky130_fd_sc_hd__o221ai_4 _08491_ (.A1(_02993_),
    .A2(_03079_),
    .B1(_03081_),
    .B2(_05576_),
    .C1(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__nor4_1 _08492_ (.A(_05590_),
    .B(_05748_),
    .C(_02967_),
    .D(_03079_),
    .Y(_03084_));
 sky130_fd_sc_hd__nor2_1 _08493_ (.A(_05572_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__mux2i_2 _08494_ (.A0(_03085_),
    .A1(_05572_),
    .S(_03083_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand3_1 _08495_ (.A(_05572_),
    .B(_02898_),
    .C(_03084_),
    .Y(_03087_));
 sky130_fd_sc_hd__o311ai_4 _08496_ (.A1(_05572_),
    .A2(_02898_),
    .A3(_03083_),
    .B1(_03086_),
    .C1(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor4_1 _08497_ (.A(_05528_),
    .B(_05774_),
    .C(_05778_),
    .D(_05787_),
    .Y(_03089_));
 sky130_fd_sc_hd__or4_1 _08498_ (.A(_05528_),
    .B(_05774_),
    .C(_05778_),
    .D(_05787_),
    .X(_03090_));
 sky130_fd_sc_hd__a21oi_1 _08499_ (.A1(_05775_),
    .A2(_03020_),
    .B1(_05779_),
    .Y(_03091_));
 sky130_fd_sc_hd__nor2_1 _08500_ (.A(_05787_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__o21bai_1 _08501_ (.A1(_05788_),
    .A2(_03092_),
    .B1_N(_05528_),
    .Y(_03093_));
 sky130_fd_sc_hd__inv_1 _08502_ (.A(_05529_),
    .Y(_03094_));
 sky130_fd_sc_hd__o211ai_1 _08503_ (.A1(_02999_),
    .A2(_03090_),
    .B1(_03093_),
    .C1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a31oi_2 _08504_ (.A1(_02906_),
    .A2(_03000_),
    .A3(_03089_),
    .B1(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__xor2_2 _08505_ (.A(_05791_),
    .B(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a22oi_4 _08506_ (.A1(_02679_),
    .A2(_03088_),
    .B1(_03097_),
    .B2(_02483_),
    .Y(_03098_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_343 ();
 sky130_fd_sc_hd__and3_4 _08508_ (.A(_02586_),
    .B(\CPU_dmem_rd_data_a5[28] ),
    .C(_01035_),
    .X(_03100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_342 ();
 sky130_fd_sc_hd__and3_1 _08510_ (.A(net1748),
    .B(_02586_),
    .C(_02596_),
    .X(_03102_));
 sky130_fd_sc_hd__a21oi_1 _08511_ (.A1(_02580_),
    .A2(_03100_),
    .B1(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__o21ai_0 _08512_ (.A1(_02582_),
    .A2(_03098_),
    .B1(_03103_),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_8 _08513_ (.A(\CPU_dmem_rd_data_a5[29] ),
    .B(_01036_),
    .Y(_03104_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_341 ();
 sky130_fd_sc_hd__clkinvlp_4 _08515_ (.A(_05795_),
    .Y(_03106_));
 sky130_fd_sc_hd__nor3_1 _08516_ (.A(_05528_),
    .B(_05770_),
    .C(_05791_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_05778_),
    .B(_05787_),
    .Y(_03108_));
 sky130_fd_sc_hd__nor2_1 _08518_ (.A(_05534_),
    .B(_05775_),
    .Y(_03109_));
 sky130_fd_sc_hd__o21ai_0 _08519_ (.A1(_05533_),
    .A2(_02976_),
    .B1(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand2b_1 _08520_ (.A_N(_05775_),
    .B(_05774_),
    .Y(_03111_));
 sky130_fd_sc_hd__inv_1 _08521_ (.A(_03065_),
    .Y(_03112_));
 sky130_fd_sc_hd__a311o_1 _08522_ (.A1(_03108_),
    .A2(_03110_),
    .A3(_03111_),
    .B1(_03112_),
    .C1(_05529_),
    .X(_03113_));
 sky130_fd_sc_hd__a21oi_1 _08523_ (.A1(_05528_),
    .A2(_03094_),
    .B1(_05791_),
    .Y(_03114_));
 sky130_fd_sc_hd__a21o_1 _08524_ (.A1(_03113_),
    .A2(_03114_),
    .B1(_05792_),
    .X(_03115_));
 sky130_fd_sc_hd__a31oi_4 _08525_ (.A1(_02917_),
    .A2(_03067_),
    .A3(_03107_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__xnor2_4 _08526_ (.A(_03106_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_340 ();
 sky130_fd_sc_hd__nor2_1 _08528_ (.A(_05572_),
    .B(_05576_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_03056_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21oi_1 _08530_ (.A1(_05576_),
    .A2(_03082_),
    .B1(_05572_),
    .Y(_03121_));
 sky130_fd_sc_hd__nor2_1 _08531_ (.A(_05573_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__a2111oi_2 _08532_ (.A1(_05582_),
    .A2(_02516_),
    .B1(_05784_),
    .C1(_05577_),
    .D1(_05573_),
    .Y(_03123_));
 sky130_fd_sc_hd__or3_1 _08533_ (.A(_05581_),
    .B(_05783_),
    .C(_03122_),
    .X(_03124_));
 sky130_fd_sc_hd__o22a_1 _08534_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03124_),
    .B2(_03013_),
    .X(_03125_));
 sky130_fd_sc_hd__inv_1 _08535_ (.A(_05567_),
    .Y(_03126_));
 sky130_fd_sc_hd__o2111a_1 _08536_ (.A1(_02967_),
    .A2(_03120_),
    .B1(_03125_),
    .C1(_03126_),
    .D1(_02679_),
    .X(_03127_));
 sky130_fd_sc_hd__nor2_1 _08537_ (.A(_05567_),
    .B(_02601_),
    .Y(_03128_));
 sky130_fd_sc_hd__o221ai_1 _08538_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03124_),
    .B2(_03013_),
    .C1(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _08539_ (.A(_05567_),
    .B(_02679_),
    .Y(_03130_));
 sky130_fd_sc_hd__o32ai_1 _08540_ (.A1(_02923_),
    .A2(_02931_),
    .A3(_03129_),
    .B1(_03130_),
    .B2(_03125_),
    .Y(_03131_));
 sky130_fd_sc_hd__and2_0 _08541_ (.A(_03056_),
    .B(_03119_),
    .X(_03132_));
 sky130_fd_sc_hd__nor2_1 _08542_ (.A(_03126_),
    .B(_02967_),
    .Y(_03133_));
 sky130_fd_sc_hd__o2111ai_1 _08543_ (.A1(_02923_),
    .A2(_02931_),
    .B1(_03132_),
    .C1(_03133_),
    .D1(_02679_),
    .Y(_03134_));
 sky130_fd_sc_hd__or3b_4 _08544_ (.A(_03127_),
    .B(_03131_),
    .C_N(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_338 ();
 sky130_fd_sc_hd__a2111oi_0 _08547_ (.A1(net98),
    .A2(_03117_),
    .B1(_02596_),
    .C1(_01035_),
    .D1(_03135_),
    .Y(_03138_));
 sky130_fd_sc_hd__nor2_1 _08548_ (.A(net1562),
    .B(_02580_),
    .Y(_03139_));
 sky130_fd_sc_hd__a2111oi_0 _08549_ (.A1(_02580_),
    .A2(_03104_),
    .B1(_03138_),
    .C1(_03139_),
    .D1(net108),
    .Y(_00565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_336 ();
 sky130_fd_sc_hd__xnor2_1 _08552_ (.A(_05641_),
    .B(_05513_),
    .Y(_03142_));
 sky130_fd_sc_hd__xnor2_1 _08553_ (.A(_05517_),
    .B(_05645_),
    .Y(_03143_));
 sky130_fd_sc_hd__o22ai_4 _08554_ (.A1(_02601_),
    .A2(_03142_),
    .B1(_03143_),
    .B2(_02632_),
    .Y(\CPU_result_a3[2] ));
 sky130_fd_sc_hd__mux2i_4 _08555_ (.A0(\CPU_dmem_rd_data_a5[2] ),
    .A1(\CPU_result_a3[2] ),
    .S(_01036_),
    .Y(_03144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_335 ();
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(_02596_),
    .B(_03144_),
    .Y(_03146_));
 sky130_fd_sc_hd__a21oi_1 _08558_ (.A1(net1621),
    .A2(_02596_),
    .B1(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__nor2_1 _08559_ (.A(net110),
    .B(_03147_),
    .Y(_00566_));
 sky130_fd_sc_hd__nor2_1 _08560_ (.A(_05567_),
    .B(_05766_),
    .Y(_03148_));
 sky130_fd_sc_hd__nand3_1 _08561_ (.A(_03043_),
    .B(_02516_),
    .C(_03046_),
    .Y(_03149_));
 sky130_fd_sc_hd__a211oi_1 _08562_ (.A1(_03123_),
    .A2(_03149_),
    .B1(_05567_),
    .C1(_03122_),
    .Y(_03150_));
 sky130_fd_sc_hd__a311oi_1 _08563_ (.A1(_02946_),
    .A2(_03132_),
    .A3(_03148_),
    .B1(_03150_),
    .C1(_05568_),
    .Y(_03151_));
 sky130_fd_sc_hd__xor2_1 _08564_ (.A(_05800_),
    .B(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__nor3_1 _08565_ (.A(_05528_),
    .B(_05791_),
    .C(_05795_),
    .Y(_03153_));
 sky130_fd_sc_hd__nor3_1 _08566_ (.A(_05528_),
    .B(_05778_),
    .C(_05787_),
    .Y(_03154_));
 sky130_fd_sc_hd__o21ai_0 _08567_ (.A1(_05528_),
    .A2(_03065_),
    .B1(_03094_),
    .Y(_03155_));
 sky130_fd_sc_hd__a21oi_1 _08568_ (.A1(_03039_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__a21oi_1 _08569_ (.A1(_05792_),
    .A2(_03106_),
    .B1(_05796_),
    .Y(_03157_));
 sky130_fd_sc_hd__o31ai_1 _08570_ (.A1(_05791_),
    .A2(_05795_),
    .A3(_03156_),
    .B1(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__a41oi_2 _08571_ (.A1(_02957_),
    .A2(_03024_),
    .A3(_03108_),
    .A4(_03153_),
    .B1(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__xor2_1 _08572_ (.A(_05804_),
    .B(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__a22oi_4 _08573_ (.A1(_02679_),
    .A2(_03152_),
    .B1(_03160_),
    .B2(_02483_),
    .Y(_03161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_334 ();
 sky130_fd_sc_hd__and3_4 _08575_ (.A(_02586_),
    .B(\CPU_dmem_rd_data_a5[30] ),
    .C(_01035_),
    .X(_03163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_333 ();
 sky130_fd_sc_hd__and3_1 _08577_ (.A(net1819),
    .B(_02586_),
    .C(_02596_),
    .X(_03165_));
 sky130_fd_sc_hd__a21oi_1 _08578_ (.A1(_02580_),
    .A2(_03163_),
    .B1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__o21ai_0 _08579_ (.A1(_02582_),
    .A2(_03161_),
    .B1(_03166_),
    .Y(_00567_));
 sky130_fd_sc_hd__nor4_1 _08580_ (.A(_05567_),
    .B(_05572_),
    .C(_05576_),
    .D(_05800_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand3_1 _08581_ (.A(_05633_),
    .B(_02679_),
    .C(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__o21bai_1 _08582_ (.A1(_05572_),
    .A2(_03082_),
    .B1_N(_05573_),
    .Y(_03169_));
 sky130_fd_sc_hd__a21oi_1 _08583_ (.A1(_03126_),
    .A2(_03169_),
    .B1(_05568_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21bai_1 _08584_ (.A1(_05800_),
    .A2(_03170_),
    .B1_N(_05801_),
    .Y(_03171_));
 sky130_fd_sc_hd__or4b_1 _08585_ (.A(_05633_),
    .B(_03171_),
    .C(_02601_),
    .D_N(_03061_),
    .X(_03172_));
 sky130_fd_sc_hd__nand2_1 _08586_ (.A(_02971_),
    .B(_03056_),
    .Y(_03173_));
 sky130_fd_sc_hd__mux2i_2 _08587_ (.A0(_03168_),
    .A1(_03172_),
    .S(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__o21bai_1 _08588_ (.A1(_03094_),
    .A2(_05791_),
    .B1_N(_05792_),
    .Y(_03175_));
 sky130_fd_sc_hd__a221oi_1 _08589_ (.A1(_03066_),
    .A2(_03153_),
    .B1(_03175_),
    .B2(_03106_),
    .C1(_05796_),
    .Y(_03176_));
 sky130_fd_sc_hd__o21bai_2 _08590_ (.A1(_05804_),
    .A2(_03176_),
    .B1_N(_05805_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand2_1 _08591_ (.A(_03067_),
    .B(_03153_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_1 _08592_ (.A(_05804_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand3_1 _08593_ (.A(_05525_),
    .B(_02483_),
    .C(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__a21oi_1 _08594_ (.A1(_02978_),
    .A2(_02980_),
    .B1(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__nor4_1 _08595_ (.A(_05525_),
    .B(_02632_),
    .C(_03177_),
    .D(_03179_),
    .Y(_03182_));
 sky130_fd_sc_hd__a311o_1 _08596_ (.A1(_05525_),
    .A2(_02483_),
    .A3(_03177_),
    .B1(_03181_),
    .C1(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__nor3_1 _08597_ (.A(_05633_),
    .B(_02601_),
    .C(_03167_),
    .Y(_03184_));
 sky130_fd_sc_hd__and2_0 _08598_ (.A(_05633_),
    .B(_02679_),
    .X(_03185_));
 sky130_fd_sc_hd__mux2i_1 _08599_ (.A0(_03184_),
    .A1(_03185_),
    .S(_03171_),
    .Y(_03186_));
 sky130_fd_sc_hd__o21a_1 _08600_ (.A1(_03061_),
    .A2(_03168_),
    .B1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o41ai_2 _08601_ (.A1(_05525_),
    .A2(_02632_),
    .A3(_02981_),
    .A4(_03177_),
    .B1(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__nor3_4 _08602_ (.A(_03174_),
    .B(_03183_),
    .C(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_332 ();
 sky130_fd_sc_hd__and3_4 _08604_ (.A(net97),
    .B(\CPU_dmem_rd_data_a5[31] ),
    .C(_01035_),
    .X(_03191_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_331 ();
 sky130_fd_sc_hd__and3_1 _08606_ (.A(net1814),
    .B(net97),
    .C(_02596_),
    .X(_03193_));
 sky130_fd_sc_hd__a21oi_1 _08607_ (.A1(_02580_),
    .A2(_03191_),
    .B1(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__o21ai_0 _08608_ (.A1(_02582_),
    .A2(_03189_),
    .B1(_03194_),
    .Y(_00568_));
 sky130_fd_sc_hd__o21bai_1 _08609_ (.A1(_05563_),
    .A2(_02647_),
    .B1_N(_05645_),
    .Y(_03195_));
 sky130_fd_sc_hd__nand2b_1 _08610_ (.A_N(_05646_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xor2_1 _08611_ (.A(_05558_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nor2_1 _08612_ (.A(_05625_),
    .B(_02667_),
    .Y(_03198_));
 sky130_fd_sc_hd__o21bai_1 _08613_ (.A1(_05641_),
    .A2(_03198_),
    .B1_N(_05642_),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_1 _08614_ (.A(_02669_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o22ai_4 _08615_ (.A1(_02632_),
    .A2(_03197_),
    .B1(_03200_),
    .B2(_02601_),
    .Y(\CPU_result_a3[3] ));
 sky130_fd_sc_hd__mux2i_4 _08616_ (.A0(\CPU_dmem_rd_data_a5[3] ),
    .A1(\CPU_result_a3[3] ),
    .S(_01036_),
    .Y(_03201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_330 ();
 sky130_fd_sc_hd__nand2_1 _08618_ (.A(net1460),
    .B(_02596_),
    .Y(_03203_));
 sky130_fd_sc_hd__o211ai_1 _08619_ (.A1(_02596_),
    .A2(_03201_),
    .B1(_03203_),
    .C1(net96),
    .Y(_00569_));
 sky130_fd_sc_hd__nor2_1 _08620_ (.A(_05558_),
    .B(_02622_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _08621_ (.A(_05559_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__xnor2_1 _08622_ (.A(_05654_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__xnor2_1 _08623_ (.A(_05650_),
    .B(_02606_),
    .Y(_03207_));
 sky130_fd_sc_hd__o22ai_4 _08624_ (.A1(_02632_),
    .A2(_03206_),
    .B1(_03207_),
    .B2(_02601_),
    .Y(\CPU_result_a3[4] ));
 sky130_fd_sc_hd__nand2_1 _08625_ (.A(_01036_),
    .B(\CPU_result_a3[4] ),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_2 _08626_ (.A(net1453),
    .B(_01035_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_8 _08627_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _08628_ (.A(_02580_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_1 _08629_ (.A(net1227),
    .B(_02596_),
    .Y(_03212_));
 sky130_fd_sc_hd__a21oi_1 _08630_ (.A1(_03211_),
    .A2(_03212_),
    .B1(net110),
    .Y(_00570_));
 sky130_fd_sc_hd__o21ai_0 _08631_ (.A1(_05621_),
    .A2(_02670_),
    .B1(_02666_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand2b_1 _08632_ (.A_N(_05651_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__xnor2_1 _08633_ (.A(_05659_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__xnor2_1 _08634_ (.A(_05663_),
    .B(_02818_),
    .Y(_03216_));
 sky130_fd_sc_hd__a22oi_4 _08635_ (.A1(_02679_),
    .A2(_03215_),
    .B1(_03216_),
    .B2(_02483_),
    .Y(_03217_));
 sky130_fd_sc_hd__nor2_1 _08636_ (.A(\CPU_dmem_rd_data_a5[5] ),
    .B(_01036_),
    .Y(_03218_));
 sky130_fd_sc_hd__a21oi_4 _08637_ (.A1(_01036_),
    .A2(_03217_),
    .B1(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _08638_ (.A(_02580_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_1 _08639_ (.A(net1224),
    .B(_02596_),
    .Y(_03221_));
 sky130_fd_sc_hd__a21oi_1 _08640_ (.A1(_03220_),
    .A2(_03221_),
    .B1(CPU_reset_a3),
    .Y(_00571_));
 sky130_fd_sc_hd__xnor2_1 _08641_ (.A(_05668_),
    .B(_02609_),
    .Y(_03222_));
 sky130_fd_sc_hd__nand2_1 _08642_ (.A(_02623_),
    .B(_02627_),
    .Y(_03223_));
 sky130_fd_sc_hd__xnor2_1 _08643_ (.A(_05672_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a22oi_4 _08644_ (.A1(_02679_),
    .A2(_03222_),
    .B1(_03224_),
    .B2(_02483_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _08645_ (.A(\CPU_dmem_rd_data_a5[6] ),
    .B(_01035_),
    .Y(_03226_));
 sky130_fd_sc_hd__o21ai_4 _08646_ (.A1(_01035_),
    .A2(_03225_),
    .B1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(_02580_),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _08648_ (.A(net1151),
    .B(_02596_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21oi_1 _08649_ (.A1(_03228_),
    .A2(_03229_),
    .B1(net109),
    .Y(_00572_));
 sky130_fd_sc_hd__a21oi_1 _08650_ (.A1(_02624_),
    .A2(_02818_),
    .B1(_05664_),
    .Y(_03230_));
 sky130_fd_sc_hd__o21bai_1 _08651_ (.A1(_05672_),
    .A2(_03230_),
    .B1_N(_05673_),
    .Y(_03231_));
 sky130_fd_sc_hd__xnor2_2 _08652_ (.A(_01080_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(_02665_),
    .B(_02673_),
    .Y(_03233_));
 sky130_fd_sc_hd__xor2_1 _08654_ (.A(_05616_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__o22ai_4 _08655_ (.A1(_02632_),
    .A2(_03232_),
    .B1(_03234_),
    .B2(_02601_),
    .Y(_03235_));
 sky130_fd_sc_hd__nor2_8 _08656_ (.A(_01035_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_329 ();
 sky130_fd_sc_hd__o21ai_4 _08658_ (.A1(\CPU_dmem_rd_data_a5[7] ),
    .A2(_01036_),
    .B1(net97),
    .Y(_03238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_327 ();
 sky130_fd_sc_hd__nand3_1 _08661_ (.A(net1613),
    .B(net96),
    .C(_02596_),
    .Y(_03241_));
 sky130_fd_sc_hd__o31ai_1 _08662_ (.A1(_02596_),
    .A2(_03236_),
    .A3(_03238_),
    .B1(_03241_),
    .Y(_00573_));
 sky130_fd_sc_hd__a31oi_1 _08663_ (.A1(_02689_),
    .A2(_02691_),
    .A3(_02692_),
    .B1(_05616_),
    .Y(_03242_));
 sky130_fd_sc_hd__nor2_1 _08664_ (.A(_05617_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__xnor2_1 _08665_ (.A(_05677_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__a211o_1 _08666_ (.A1(_02623_),
    .A2(_02627_),
    .B1(_05553_),
    .C1(_05672_),
    .X(_03245_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_02618_),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__xnor2_1 _08668_ (.A(_02655_),
    .B(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__o22ai_4 _08669_ (.A1(_02601_),
    .A2(_03244_),
    .B1(_03247_),
    .B2(_02632_),
    .Y(_03248_));
 sky130_fd_sc_hd__nor2_1 _08670_ (.A(_01035_),
    .B(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__nor2_1 _08671_ (.A(\CPU_dmem_rd_data_a5[8] ),
    .B(_01036_),
    .Y(_03250_));
 sky130_fd_sc_hd__or3_4 _08672_ (.A(CPU_reset_a3),
    .B(_03249_),
    .C(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_326 ();
 sky130_fd_sc_hd__nand3_1 _08674_ (.A(net1421),
    .B(net96),
    .C(_02596_),
    .Y(_03253_));
 sky130_fd_sc_hd__o21ai_0 _08675_ (.A1(_02596_),
    .A2(_03251_),
    .B1(_03253_),
    .Y(_00574_));
 sky130_fd_sc_hd__nor2_1 _08676_ (.A(_02663_),
    .B(_02674_),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _08677_ (.A(_05686_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__nor2_1 _08678_ (.A(_02652_),
    .B(_02657_),
    .Y(_03256_));
 sky130_fd_sc_hd__xnor2_2 _08679_ (.A(_05690_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__o22ai_4 _08680_ (.A1(_02601_),
    .A2(_03255_),
    .B1(_03257_),
    .B2(_02632_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_8 _08681_ (.A(_01035_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_325 ();
 sky130_fd_sc_hd__o21ai_4 _08683_ (.A1(\CPU_dmem_rd_data_a5[9] ),
    .A2(_01036_),
    .B1(net96),
    .Y(_03261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_324 ();
 sky130_fd_sc_hd__nand3_1 _08685_ (.A(net1332),
    .B(net96),
    .C(_02596_),
    .Y(_03263_));
 sky130_fd_sc_hd__o31ai_1 _08686_ (.A1(_02596_),
    .A2(_03259_),
    .A3(_03261_),
    .B1(_03263_),
    .Y(_00575_));
 sky130_fd_sc_hd__nor2_1 _08687_ (.A(\CPU_dmem_rd_data_a5[0] ),
    .B(_01036_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21o_2 _08688_ (.A1(_01036_),
    .A2(_02560_),
    .B1(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__nand3_1 _08689_ (.A(\CPU_rd_a3[0] ),
    .B(\CPU_rd_a3[1] ),
    .C(_01036_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand3_1 _08690_ (.A(\CPU_rd_a5[0] ),
    .B(\CPU_rd_a5[1] ),
    .C(_01035_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_4 _08691_ (.A(_03266_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__and2_4 _08692_ (.A(_02574_),
    .B(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__nand2_8 _08693_ (.A(_02592_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_320 ();
 sky130_fd_sc_hd__a21oi_1 _08698_ (.A1(net1652),
    .A2(_03270_),
    .B1(CPU_reset_a3),
    .Y(_03275_));
 sky130_fd_sc_hd__o21ai_0 _08699_ (.A1(_03265_),
    .A2(_03270_),
    .B1(_03275_),
    .Y(_00576_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_319 ();
 sky130_fd_sc_hd__nand2_4 _08701_ (.A(_02574_),
    .B(_03268_),
    .Y(_03277_));
 sky130_fd_sc_hd__nor2_8 _08702_ (.A(_02567_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_318 ();
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(_02636_),
    .B(_03278_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(net1306),
    .B(_03270_),
    .Y(_03281_));
 sky130_fd_sc_hd__a21oi_1 _08706_ (.A1(_03280_),
    .A2(_03281_),
    .B1(net108),
    .Y(_00577_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_317 ();
 sky130_fd_sc_hd__nand2_1 _08708_ (.A(net1134),
    .B(_03270_),
    .Y(_03283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_316 ();
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_02683_),
    .B(_03278_),
    .Y(_03285_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_315 ();
 sky130_fd_sc_hd__a21oi_1 _08712_ (.A1(_03283_),
    .A2(_03285_),
    .B1(net109),
    .Y(_00578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_313 ();
 sky130_fd_sc_hd__nand3_1 _08715_ (.A(net1469),
    .B(net96),
    .C(_03270_),
    .Y(_03289_));
 sky130_fd_sc_hd__o21ai_0 _08716_ (.A1(_02713_),
    .A2(_03270_),
    .B1(_03289_),
    .Y(_00579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_312 ();
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_02748_),
    .B(_03278_),
    .Y(_03291_));
 sky130_fd_sc_hd__nand2_1 _08719_ (.A(net1092),
    .B(_03270_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _08720_ (.A1(_03291_),
    .A2(_03292_),
    .B1(net109),
    .Y(_00580_));
 sky130_fd_sc_hd__nand3_1 _08721_ (.A(net1394),
    .B(net97),
    .C(_03270_),
    .Y(_03293_));
 sky130_fd_sc_hd__o21ai_0 _08722_ (.A1(_02766_),
    .A2(_03270_),
    .B1(_03293_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand3_1 _08723_ (.A(net1628),
    .B(net97),
    .C(_03270_),
    .Y(_03294_));
 sky130_fd_sc_hd__o21ai_0 _08724_ (.A1(_02784_),
    .A2(_03270_),
    .B1(_03294_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand3_1 _08725_ (.A(net1454),
    .B(net97),
    .C(_03270_),
    .Y(_03295_));
 sky130_fd_sc_hd__o21ai_0 _08726_ (.A1(_02809_),
    .A2(_03270_),
    .B1(_03295_),
    .Y(_00583_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_311 ();
 sky130_fd_sc_hd__nand2_8 _08728_ (.A(_02581_),
    .B(_03278_),
    .Y(_03297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_310 ();
 sky130_fd_sc_hd__nand3_1 _08730_ (.A(net1531),
    .B(net97),
    .C(_03270_),
    .Y(_03299_));
 sky130_fd_sc_hd__o221ai_1 _08731_ (.A1(_02834_),
    .A2(_03270_),
    .B1(_03297_),
    .B2(_02832_),
    .C1(_03299_),
    .Y(_00584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_308 ();
 sky130_fd_sc_hd__and3_1 _08734_ (.A(net1727),
    .B(_02586_),
    .C(_03270_),
    .X(_03302_));
 sky130_fd_sc_hd__a31o_1 _08735_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03278_),
    .B1(_03302_),
    .X(_00585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_307 ();
 sky130_fd_sc_hd__and3_1 _08737_ (.A(net1742),
    .B(net97),
    .C(_03270_),
    .X(_03304_));
 sky130_fd_sc_hd__a21oi_1 _08738_ (.A1(_02884_),
    .A2(_03278_),
    .B1(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__o21ai_0 _08739_ (.A1(_02882_),
    .A2(_03297_),
    .B1(_03305_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(net1488),
    .B(_03270_),
    .Y(_03306_));
 sky130_fd_sc_hd__o211ai_1 _08741_ (.A1(_02889_),
    .A2(_03270_),
    .B1(_03306_),
    .C1(_02586_),
    .Y(_00587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_306 ();
 sky130_fd_sc_hd__nand3_1 _08743_ (.A(net1629),
    .B(net97),
    .C(_03270_),
    .Y(_03308_));
 sky130_fd_sc_hd__o221ai_1 _08744_ (.A1(_02909_),
    .A2(_03270_),
    .B1(_03297_),
    .B2(_02908_),
    .C1(_03308_),
    .Y(_00588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_305 ();
 sky130_fd_sc_hd__nand3_1 _08746_ (.A(net1580),
    .B(_02586_),
    .C(_03270_),
    .Y(_03310_));
 sky130_fd_sc_hd__o221ai_1 _08747_ (.A1(_02936_),
    .A2(_03270_),
    .B1(_03297_),
    .B2(_02934_),
    .C1(_03310_),
    .Y(_00589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_304 ();
 sky130_fd_sc_hd__and3_1 _08749_ (.A(net1783),
    .B(_02586_),
    .C(_03270_),
    .X(_03312_));
 sky130_fd_sc_hd__a21oi_1 _08750_ (.A1(_02961_),
    .A2(_03278_),
    .B1(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__o21ai_0 _08751_ (.A1(_02959_),
    .A2(_03297_),
    .B1(_03313_),
    .Y(_00590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_303 ();
 sky130_fd_sc_hd__nand3_1 _08753_ (.A(net1589),
    .B(net97),
    .C(_03270_),
    .Y(_03315_));
 sky130_fd_sc_hd__o221ai_1 _08754_ (.A1(_02984_),
    .A2(_03270_),
    .B1(_03297_),
    .B2(_02983_),
    .C1(_03315_),
    .Y(_00591_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_302 ();
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_03009_),
    .B(_03278_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_1 _08757_ (.A(net1241),
    .B(_03270_),
    .Y(_03318_));
 sky130_fd_sc_hd__a21oi_1 _08758_ (.A1(_03317_),
    .A2(_03318_),
    .B1(net109),
    .Y(_00592_));
 sky130_fd_sc_hd__nor2_1 _08759_ (.A(_01035_),
    .B(_03270_),
    .Y(_03319_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_301 ();
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_03031_),
    .B(_03278_),
    .Y(_03321_));
 sky130_fd_sc_hd__o21ai_0 _08762_ (.A1(net1714),
    .A2(_03278_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__a311oi_1 _08763_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03319_),
    .B1(_03322_),
    .C1(net108),
    .Y(_00593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_300 ();
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_03053_),
    .B(_03278_),
    .Y(_03324_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(net1337),
    .B(_03270_),
    .Y(_03325_));
 sky130_fd_sc_hd__a21oi_1 _08767_ (.A1(_03324_),
    .A2(_03325_),
    .B1(net109),
    .Y(_00594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_299 ();
 sky130_fd_sc_hd__nand3_1 _08769_ (.A(net1484),
    .B(_02586_),
    .C(_03270_),
    .Y(_03327_));
 sky130_fd_sc_hd__o221ai_1 _08770_ (.A1(_03076_),
    .A2(_03270_),
    .B1(_03297_),
    .B2(_03074_),
    .C1(_03327_),
    .Y(_00595_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_298 ();
 sky130_fd_sc_hd__and3_1 _08772_ (.A(net1815),
    .B(_02586_),
    .C(_03270_),
    .X(_03329_));
 sky130_fd_sc_hd__a21oi_1 _08773_ (.A1(_03100_),
    .A2(_03278_),
    .B1(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__o21ai_0 _08774_ (.A1(_03098_),
    .A2(_03297_),
    .B1(_03330_),
    .Y(_00596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_296 ();
 sky130_fd_sc_hd__a2111oi_0 _08777_ (.A1(net98),
    .A2(_03117_),
    .B1(_03270_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03333_));
 sky130_fd_sc_hd__nor2_1 _08778_ (.A(net1614),
    .B(_03278_),
    .Y(_03334_));
 sky130_fd_sc_hd__a2111oi_0 _08779_ (.A1(_03104_),
    .A2(_03278_),
    .B1(_03333_),
    .C1(_03334_),
    .D1(net108),
    .Y(_00597_));
 sky130_fd_sc_hd__nor2_1 _08780_ (.A(_03144_),
    .B(_03270_),
    .Y(_03335_));
 sky130_fd_sc_hd__a21oi_1 _08781_ (.A1(net1662),
    .A2(_03270_),
    .B1(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__nor2_1 _08782_ (.A(net110),
    .B(_03336_),
    .Y(_00598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_294 ();
 sky130_fd_sc_hd__and3_1 _08785_ (.A(net1804),
    .B(_02586_),
    .C(_03270_),
    .X(_03339_));
 sky130_fd_sc_hd__a21oi_1 _08786_ (.A1(_03163_),
    .A2(_03278_),
    .B1(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__o21ai_0 _08787_ (.A1(_03161_),
    .A2(_03297_),
    .B1(_03340_),
    .Y(_00599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_293 ();
 sky130_fd_sc_hd__and3_1 _08789_ (.A(net1808),
    .B(net97),
    .C(_03270_),
    .X(_03342_));
 sky130_fd_sc_hd__a21oi_1 _08790_ (.A1(_03191_),
    .A2(_03278_),
    .B1(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21ai_0 _08791_ (.A1(_03189_),
    .A2(_03297_),
    .B1(_03343_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(net1507),
    .B(_03270_),
    .Y(_03344_));
 sky130_fd_sc_hd__o211ai_1 _08793_ (.A1(_03201_),
    .A2(_03270_),
    .B1(_03344_),
    .C1(net96),
    .Y(_00601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_292 ();
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(_03210_),
    .B(_03278_),
    .Y(_03346_));
 sky130_fd_sc_hd__nand2_1 _08796_ (.A(net1217),
    .B(_03270_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_1 _08797_ (.A1(_03346_),
    .A2(_03347_),
    .B1(net110),
    .Y(_00602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_291 ();
 sky130_fd_sc_hd__nand2_1 _08799_ (.A(_03219_),
    .B(_03278_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(net1283),
    .B(_03270_),
    .Y(_03350_));
 sky130_fd_sc_hd__a21oi_1 _08801_ (.A1(_03349_),
    .A2(_03350_),
    .B1(net110),
    .Y(_00603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_290 ();
 sky130_fd_sc_hd__nand2_1 _08803_ (.A(_03227_),
    .B(_03278_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand2_1 _08804_ (.A(net1225),
    .B(_03270_),
    .Y(_03353_));
 sky130_fd_sc_hd__a21oi_1 _08805_ (.A1(_03352_),
    .A2(_03353_),
    .B1(net110),
    .Y(_00604_));
 sky130_fd_sc_hd__nand3_1 _08806_ (.A(net1416),
    .B(net96),
    .C(_03270_),
    .Y(_03354_));
 sky130_fd_sc_hd__o31ai_1 _08807_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03270_),
    .B1(_03354_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand3_1 _08808_ (.A(net1437),
    .B(net96),
    .C(_03270_),
    .Y(_03355_));
 sky130_fd_sc_hd__o21ai_0 _08809_ (.A1(_03251_),
    .A2(_03270_),
    .B1(_03355_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand3_1 _08810_ (.A(net1431),
    .B(net96),
    .C(_03270_),
    .Y(_03356_));
 sky130_fd_sc_hd__o31ai_1 _08811_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03270_),
    .B1(_03356_),
    .Y(_00607_));
 sky130_fd_sc_hd__and3_1 _08812_ (.A(\CPU_rd_a5[2] ),
    .B(\CPU_rd_a5[3] ),
    .C(_01035_),
    .X(_03357_));
 sky130_fd_sc_hd__a31oi_4 _08813_ (.A1(\CPU_rd_a3[2] ),
    .A2(\CPU_rd_a3[3] ),
    .A3(_01036_),
    .B1(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nor3_1 _08814_ (.A(\CPU_rd_a5[0] ),
    .B(\CPU_rd_a5[1] ),
    .C(_01036_),
    .Y(_03359_));
 sky130_fd_sc_hd__a21o_1 _08815_ (.A1(_01036_),
    .A2(_02570_),
    .B1(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__nand2_4 _08816_ (.A(_02574_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__nor2_8 _08817_ (.A(_03358_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_8 _08818_ (.A(_02581_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_287 ();
 sky130_fd_sc_hd__a31o_4 _08822_ (.A1(\CPU_rd_a3[2] ),
    .A2(\CPU_rd_a3[3] ),
    .A3(_01036_),
    .B1(_03357_),
    .X(_03367_));
 sky130_fd_sc_hd__and2_4 _08823_ (.A(_02574_),
    .B(_03360_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_8 _08824_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_286 ();
 sky130_fd_sc_hd__and3_1 _08826_ (.A(net1807),
    .B(net97),
    .C(_03369_),
    .X(_03371_));
 sky130_fd_sc_hd__a21oi_1 _08827_ (.A1(_02588_),
    .A2(_03362_),
    .B1(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__o21ai_0 _08828_ (.A1(_02560_),
    .A2(_03363_),
    .B1(_03372_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _08829_ (.A(_02636_),
    .B(_03362_),
    .Y(_03373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_285 ();
 sky130_fd_sc_hd__nand2_1 _08831_ (.A(net1236),
    .B(_03369_),
    .Y(_03375_));
 sky130_fd_sc_hd__a21oi_1 _08832_ (.A1(_03373_),
    .A2(_03375_),
    .B1(net108),
    .Y(_00609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_284 ();
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(net1340),
    .B(_03369_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_02683_),
    .B(_03362_),
    .Y(_03378_));
 sky130_fd_sc_hd__a21oi_1 _08836_ (.A1(_03377_),
    .A2(_03378_),
    .B1(net109),
    .Y(_00610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_282 ();
 sky130_fd_sc_hd__nand3_1 _08839_ (.A(net1481),
    .B(net96),
    .C(_03369_),
    .Y(_03381_));
 sky130_fd_sc_hd__o21ai_0 _08840_ (.A1(_02713_),
    .A2(_03369_),
    .B1(_03381_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_02748_),
    .B(_03362_),
    .Y(_03382_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(net1234),
    .B(_03369_),
    .Y(_03383_));
 sky130_fd_sc_hd__a21oi_1 _08843_ (.A1(_03382_),
    .A2(_03383_),
    .B1(net109),
    .Y(_00612_));
 sky130_fd_sc_hd__nand3_1 _08844_ (.A(net1426),
    .B(net97),
    .C(_03369_),
    .Y(_03384_));
 sky130_fd_sc_hd__o21ai_0 _08845_ (.A1(_02766_),
    .A2(_03369_),
    .B1(_03384_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand3_1 _08846_ (.A(net1367),
    .B(net97),
    .C(_03369_),
    .Y(_03385_));
 sky130_fd_sc_hd__o21ai_0 _08847_ (.A1(_02784_),
    .A2(_03369_),
    .B1(_03385_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand3_1 _08848_ (.A(net1403),
    .B(net97),
    .C(_03369_),
    .Y(_03386_));
 sky130_fd_sc_hd__o21ai_0 _08849_ (.A1(_02809_),
    .A2(_03369_),
    .B1(_03386_),
    .Y(_00615_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_281 ();
 sky130_fd_sc_hd__nand3_1 _08851_ (.A(net1566),
    .B(net97),
    .C(_03369_),
    .Y(_03388_));
 sky130_fd_sc_hd__o221ai_1 _08852_ (.A1(_02834_),
    .A2(_03369_),
    .B1(_03363_),
    .B2(_02832_),
    .C1(_03388_),
    .Y(_00616_));
 sky130_fd_sc_hd__and3_1 _08853_ (.A(net1710),
    .B(_02586_),
    .C(_03369_),
    .X(_03389_));
 sky130_fd_sc_hd__a31o_1 _08854_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03362_),
    .B1(_03389_),
    .X(_00617_));
 sky130_fd_sc_hd__and3_1 _08855_ (.A(net1743),
    .B(net97),
    .C(_03369_),
    .X(_03390_));
 sky130_fd_sc_hd__a21oi_1 _08856_ (.A1(_02884_),
    .A2(_03362_),
    .B1(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__o21ai_0 _08857_ (.A1(_02882_),
    .A2(_03363_),
    .B1(_03391_),
    .Y(_00618_));
 sky130_fd_sc_hd__nor2_1 _08858_ (.A(_02889_),
    .B(_03369_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21oi_1 _08859_ (.A1(net1491),
    .A2(_03369_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_1 _08860_ (.A(CPU_reset_a3),
    .B(_03393_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand3_1 _08861_ (.A(net1553),
    .B(net96),
    .C(_03369_),
    .Y(_03394_));
 sky130_fd_sc_hd__o221ai_1 _08862_ (.A1(_02909_),
    .A2(_03369_),
    .B1(_03363_),
    .B2(_02908_),
    .C1(_03394_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand3_1 _08863_ (.A(net1598),
    .B(net96),
    .C(_03369_),
    .Y(_03395_));
 sky130_fd_sc_hd__o221ai_1 _08864_ (.A1(_02936_),
    .A2(_03369_),
    .B1(_03363_),
    .B2(_02934_),
    .C1(_03395_),
    .Y(_00621_));
 sky130_fd_sc_hd__and3_1 _08865_ (.A(net1779),
    .B(_02586_),
    .C(_03369_),
    .X(_03396_));
 sky130_fd_sc_hd__a21oi_1 _08866_ (.A1(_02961_),
    .A2(_03362_),
    .B1(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21ai_0 _08867_ (.A1(_02959_),
    .A2(_03363_),
    .B1(_03397_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand3_1 _08868_ (.A(net1655),
    .B(net97),
    .C(_03369_),
    .Y(_03398_));
 sky130_fd_sc_hd__o221ai_1 _08869_ (.A1(_02984_),
    .A2(_03369_),
    .B1(_03363_),
    .B2(_02983_),
    .C1(_03398_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_03009_),
    .B(_03362_),
    .Y(_03399_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(net1216),
    .B(_03369_),
    .Y(_03400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_280 ();
 sky130_fd_sc_hd__a21oi_1 _08873_ (.A1(_03399_),
    .A2(_03400_),
    .B1(net109),
    .Y(_00624_));
 sky130_fd_sc_hd__nor2_1 _08874_ (.A(_01035_),
    .B(_03369_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(_03031_),
    .B(_03362_),
    .Y(_03403_));
 sky130_fd_sc_hd__o21ai_0 _08876_ (.A1(net1692),
    .A2(_03362_),
    .B1(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__a311oi_1 _08877_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03402_),
    .B1(_03404_),
    .C1(net108),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _08878_ (.A(_03053_),
    .B(_03362_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(net1201),
    .B(_03369_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21oi_1 _08880_ (.A1(_03405_),
    .A2(_03406_),
    .B1(net109),
    .Y(_00626_));
 sky130_fd_sc_hd__nand3_1 _08881_ (.A(net1623),
    .B(net97),
    .C(_03369_),
    .Y(_03407_));
 sky130_fd_sc_hd__o221ai_1 _08882_ (.A1(_03076_),
    .A2(_03369_),
    .B1(_03363_),
    .B2(_03074_),
    .C1(_03407_),
    .Y(_00627_));
 sky130_fd_sc_hd__and3_1 _08883_ (.A(net1839),
    .B(net97),
    .C(_03369_),
    .X(_03408_));
 sky130_fd_sc_hd__a21oi_1 _08884_ (.A1(_03100_),
    .A2(_03362_),
    .B1(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__o21ai_0 _08885_ (.A1(_03098_),
    .A2(_03363_),
    .B1(_03409_),
    .Y(_00628_));
 sky130_fd_sc_hd__a2111oi_0 _08886_ (.A1(net98),
    .A2(_03117_),
    .B1(_03369_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03410_));
 sky130_fd_sc_hd__nor2_1 _08887_ (.A(net1680),
    .B(_03362_),
    .Y(_03411_));
 sky130_fd_sc_hd__a2111oi_0 _08888_ (.A1(_03104_),
    .A2(_03362_),
    .B1(_03410_),
    .C1(_03411_),
    .D1(net108),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _08889_ (.A(net1461),
    .B(_03369_),
    .Y(_03412_));
 sky130_fd_sc_hd__o211ai_1 _08890_ (.A1(_03144_),
    .A2(_03369_),
    .B1(_03412_),
    .C1(net96),
    .Y(_00630_));
 sky130_fd_sc_hd__and3_1 _08891_ (.A(net1806),
    .B(_02586_),
    .C(_03369_),
    .X(_03413_));
 sky130_fd_sc_hd__a21oi_1 _08892_ (.A1(_03163_),
    .A2(_03362_),
    .B1(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_0 _08893_ (.A1(_03161_),
    .A2(_03363_),
    .B1(_03414_),
    .Y(_00631_));
 sky130_fd_sc_hd__and3_1 _08894_ (.A(net1729),
    .B(net97),
    .C(_03369_),
    .X(_03415_));
 sky130_fd_sc_hd__a21oi_1 _08895_ (.A1(_03191_),
    .A2(_03362_),
    .B1(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21ai_0 _08896_ (.A1(_03189_),
    .A2(_03363_),
    .B1(_03416_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(net1465),
    .B(_03369_),
    .Y(_03417_));
 sky130_fd_sc_hd__o211ai_1 _08898_ (.A1(_03201_),
    .A2(_03369_),
    .B1(_03417_),
    .C1(net96),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(_03210_),
    .B(_03362_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(net1285),
    .B(_03369_),
    .Y(_03419_));
 sky130_fd_sc_hd__a21oi_1 _08901_ (.A1(_03418_),
    .A2(_03419_),
    .B1(net110),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _08902_ (.A(_03219_),
    .B(_03362_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_1 _08903_ (.A(net1427),
    .B(_03369_),
    .Y(_03421_));
 sky130_fd_sc_hd__a21oi_1 _08904_ (.A1(_03420_),
    .A2(_03421_),
    .B1(CPU_reset_a3),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _08905_ (.A(_03227_),
    .B(_03362_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand2_1 _08906_ (.A(net1296),
    .B(_03369_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_1 _08907_ (.A1(_03422_),
    .A2(_03423_),
    .B1(net110),
    .Y(_00636_));
 sky130_fd_sc_hd__nand3_1 _08908_ (.A(net1368),
    .B(net96),
    .C(_03369_),
    .Y(_03424_));
 sky130_fd_sc_hd__o31ai_1 _08909_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03369_),
    .B1(_03424_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand3_1 _08910_ (.A(net1436),
    .B(net96),
    .C(_03369_),
    .Y(_03425_));
 sky130_fd_sc_hd__o21ai_0 _08911_ (.A1(_03251_),
    .A2(_03369_),
    .B1(_03425_),
    .Y(_00638_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_279 ();
 sky130_fd_sc_hd__nand3_1 _08913_ (.A(net1323),
    .B(net96),
    .C(_03369_),
    .Y(_03427_));
 sky130_fd_sc_hd__o31ai_1 _08914_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03369_),
    .B1(_03427_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2b_1 _08915_ (.A_N(\CPU_rd_a5[1] ),
    .B(\CPU_rd_a5[0] ),
    .Y(_03428_));
 sky130_fd_sc_hd__or3_1 _08916_ (.A(_02576_),
    .B(\CPU_rd_a3[1] ),
    .C(_01035_),
    .X(_03429_));
 sky130_fd_sc_hd__o21a_2 _08917_ (.A1(_01036_),
    .A2(_03428_),
    .B1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nor2_8 _08918_ (.A(_02593_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_8 _08919_ (.A(_03367_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_276 ();
 sky130_fd_sc_hd__a21oi_1 _08923_ (.A1(net1608),
    .A2(_03432_),
    .B1(net108),
    .Y(_03436_));
 sky130_fd_sc_hd__o21ai_0 _08924_ (.A1(_03265_),
    .A2(_03432_),
    .B1(_03436_),
    .Y(_00640_));
 sky130_fd_sc_hd__o21ai_4 _08925_ (.A1(_01036_),
    .A2(_03428_),
    .B1(_03429_),
    .Y(_03437_));
 sky130_fd_sc_hd__nand2_4 _08926_ (.A(_02574_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__nor2_8 _08927_ (.A(_03358_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_275 ();
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(_02636_),
    .B(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _08930_ (.A(net1089),
    .B(_03432_),
    .Y(_03442_));
 sky130_fd_sc_hd__a21oi_1 _08931_ (.A1(_03441_),
    .A2(_03442_),
    .B1(net108),
    .Y(_00641_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 ();
 sky130_fd_sc_hd__nand2_1 _08933_ (.A(net1315),
    .B(_03432_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(_02683_),
    .B(_03439_),
    .Y(_03445_));
 sky130_fd_sc_hd__a21oi_1 _08935_ (.A1(_03444_),
    .A2(_03445_),
    .B1(net109),
    .Y(_00642_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_272 ();
 sky130_fd_sc_hd__nand3_1 _08938_ (.A(net1546),
    .B(net96),
    .C(_03432_),
    .Y(_03448_));
 sky130_fd_sc_hd__o21ai_0 _08939_ (.A1(_02713_),
    .A2(_03432_),
    .B1(_03448_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _08940_ (.A(_02748_),
    .B(_03439_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _08941_ (.A(net1391),
    .B(_03432_),
    .Y(_03450_));
 sky130_fd_sc_hd__a21oi_1 _08942_ (.A1(_03449_),
    .A2(_03450_),
    .B1(net109),
    .Y(_00644_));
 sky130_fd_sc_hd__nand3_1 _08943_ (.A(net1476),
    .B(net97),
    .C(_03432_),
    .Y(_03451_));
 sky130_fd_sc_hd__o21ai_0 _08944_ (.A1(_02766_),
    .A2(_03432_),
    .B1(_03451_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand3_1 _08945_ (.A(net1496),
    .B(net97),
    .C(_03432_),
    .Y(_03452_));
 sky130_fd_sc_hd__o21ai_0 _08946_ (.A1(_02784_),
    .A2(_03432_),
    .B1(_03452_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand3_1 _08947_ (.A(net1380),
    .B(net97),
    .C(_03432_),
    .Y(_03453_));
 sky130_fd_sc_hd__o21ai_0 _08948_ (.A1(_02809_),
    .A2(_03432_),
    .B1(_03453_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_8 _08949_ (.A(_02581_),
    .B(_03439_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand3_1 _08950_ (.A(net1602),
    .B(net97),
    .C(_03432_),
    .Y(_03455_));
 sky130_fd_sc_hd__o221ai_1 _08951_ (.A1(_02834_),
    .A2(_03432_),
    .B1(_03454_),
    .B2(_02832_),
    .C1(_03455_),
    .Y(_00648_));
 sky130_fd_sc_hd__and3_1 _08952_ (.A(net1838),
    .B(_02586_),
    .C(_03432_),
    .X(_03456_));
 sky130_fd_sc_hd__a31o_1 _08953_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03439_),
    .B1(_03456_),
    .X(_00649_));
 sky130_fd_sc_hd__and3_1 _08954_ (.A(net1741),
    .B(net97),
    .C(_03432_),
    .X(_03457_));
 sky130_fd_sc_hd__a21oi_1 _08955_ (.A1(_02884_),
    .A2(_03439_),
    .B1(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__o21ai_0 _08956_ (.A1(_02882_),
    .A2(_03454_),
    .B1(_03458_),
    .Y(_00650_));
 sky130_fd_sc_hd__nor2_1 _08957_ (.A(_02889_),
    .B(_03432_),
    .Y(_03459_));
 sky130_fd_sc_hd__a21oi_1 _08958_ (.A1(net1624),
    .A2(_03432_),
    .B1(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__nor2_1 _08959_ (.A(net110),
    .B(_03460_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand3_1 _08960_ (.A(net1647),
    .B(net97),
    .C(_03432_),
    .Y(_03461_));
 sky130_fd_sc_hd__o221ai_1 _08961_ (.A1(_02909_),
    .A2(_03432_),
    .B1(_03454_),
    .B2(_02908_),
    .C1(_03461_),
    .Y(_00652_));
 sky130_fd_sc_hd__nand3_1 _08962_ (.A(net1612),
    .B(_02586_),
    .C(_03432_),
    .Y(_03462_));
 sky130_fd_sc_hd__o221ai_1 _08963_ (.A1(_02936_),
    .A2(_03432_),
    .B1(_03454_),
    .B2(_02934_),
    .C1(_03462_),
    .Y(_00653_));
 sky130_fd_sc_hd__and3_1 _08964_ (.A(net1756),
    .B(_02586_),
    .C(_03432_),
    .X(_03463_));
 sky130_fd_sc_hd__a21oi_1 _08965_ (.A1(_02961_),
    .A2(_03439_),
    .B1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__o21ai_0 _08966_ (.A1(_02959_),
    .A2(_03454_),
    .B1(_03464_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand3_1 _08967_ (.A(net1664),
    .B(_02586_),
    .C(_03432_),
    .Y(_03465_));
 sky130_fd_sc_hd__o221ai_1 _08968_ (.A1(_02984_),
    .A2(_03432_),
    .B1(_03454_),
    .B2(_02983_),
    .C1(_03465_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_03009_),
    .B(_03439_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(net1372),
    .B(_03432_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21oi_1 _08971_ (.A1(_03466_),
    .A2(_03467_),
    .B1(net109),
    .Y(_00656_));
 sky130_fd_sc_hd__nor2_1 _08972_ (.A(_01035_),
    .B(_03432_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _08973_ (.A(_03031_),
    .B(_03439_),
    .Y(_03469_));
 sky130_fd_sc_hd__o21ai_0 _08974_ (.A1(net1721),
    .A2(_03439_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__a311oi_1 _08975_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03468_),
    .B1(_03470_),
    .C1(net108),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(_03053_),
    .B(_03439_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _08977_ (.A(net1411),
    .B(_03432_),
    .Y(_03472_));
 sky130_fd_sc_hd__a21oi_1 _08978_ (.A1(_03471_),
    .A2(_03472_),
    .B1(net109),
    .Y(_00658_));
 sky130_fd_sc_hd__nand3_1 _08979_ (.A(net1601),
    .B(_02586_),
    .C(_03432_),
    .Y(_03473_));
 sky130_fd_sc_hd__o221ai_1 _08980_ (.A1(_03076_),
    .A2(_03432_),
    .B1(_03454_),
    .B2(_03074_),
    .C1(_03473_),
    .Y(_00659_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_271 ();
 sky130_fd_sc_hd__and3_1 _08982_ (.A(net1782),
    .B(net97),
    .C(_03432_),
    .X(_03475_));
 sky130_fd_sc_hd__a21oi_1 _08983_ (.A1(_03100_),
    .A2(_03439_),
    .B1(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__o21ai_0 _08984_ (.A1(_03098_),
    .A2(_03454_),
    .B1(_03476_),
    .Y(_00660_));
 sky130_fd_sc_hd__a2111oi_0 _08985_ (.A1(net98),
    .A2(_03117_),
    .B1(_03432_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03477_));
 sky130_fd_sc_hd__nor2_1 _08986_ (.A(net1535),
    .B(_03439_),
    .Y(_03478_));
 sky130_fd_sc_hd__a2111oi_0 _08987_ (.A1(_03104_),
    .A2(_03439_),
    .B1(_03477_),
    .C1(_03478_),
    .D1(net108),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(net1492),
    .B(_03432_),
    .Y(_03479_));
 sky130_fd_sc_hd__o211ai_1 _08989_ (.A1(_03144_),
    .A2(_03432_),
    .B1(_03479_),
    .C1(_02586_),
    .Y(_00662_));
 sky130_fd_sc_hd__and3_1 _08990_ (.A(net1758),
    .B(_02586_),
    .C(_03432_),
    .X(_03480_));
 sky130_fd_sc_hd__a21oi_1 _08991_ (.A1(_03163_),
    .A2(_03439_),
    .B1(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__o21ai_0 _08992_ (.A1(_03161_),
    .A2(_03454_),
    .B1(_03481_),
    .Y(_00663_));
 sky130_fd_sc_hd__and3_1 _08993_ (.A(net1843),
    .B(net97),
    .C(_03432_),
    .X(_03482_));
 sky130_fd_sc_hd__a21oi_1 _08994_ (.A1(_03191_),
    .A2(_03439_),
    .B1(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__o21ai_0 _08995_ (.A1(_03189_),
    .A2(_03454_),
    .B1(_03483_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(net1576),
    .B(_03432_),
    .Y(_03484_));
 sky130_fd_sc_hd__o211ai_1 _08997_ (.A1(_03201_),
    .A2(_03432_),
    .B1(_03484_),
    .C1(net96),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(_03210_),
    .B(_03439_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _08999_ (.A(net1197),
    .B(_03432_),
    .Y(_03486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_270 ();
 sky130_fd_sc_hd__a21oi_1 _09001_ (.A1(_03485_),
    .A2(_03486_),
    .B1(net110),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(_03219_),
    .B(_03439_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(net1334),
    .B(_03432_),
    .Y(_03489_));
 sky130_fd_sc_hd__a21oi_1 _09004_ (.A1(_03488_),
    .A2(_03489_),
    .B1(CPU_reset_a3),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_03227_),
    .B(_03439_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(net1245),
    .B(_03432_),
    .Y(_03491_));
 sky130_fd_sc_hd__a21oi_1 _09007_ (.A1(_03490_),
    .A2(_03491_),
    .B1(net109),
    .Y(_00668_));
 sky130_fd_sc_hd__nand3_1 _09008_ (.A(net1493),
    .B(net96),
    .C(_03432_),
    .Y(_03492_));
 sky130_fd_sc_hd__o31ai_1 _09009_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03432_),
    .B1(_03492_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand3_1 _09010_ (.A(net1420),
    .B(net96),
    .C(_03432_),
    .Y(_03493_));
 sky130_fd_sc_hd__o21ai_0 _09011_ (.A1(_03251_),
    .A2(_03432_),
    .B1(_03493_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand3_1 _09012_ (.A(net1443),
    .B(net96),
    .C(_03432_),
    .Y(_03494_));
 sky130_fd_sc_hd__o31ai_1 _09013_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03432_),
    .B1(_03494_),
    .Y(_00671_));
 sky130_fd_sc_hd__nor2_8 _09014_ (.A(_02579_),
    .B(_03358_),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_8 _09015_ (.A(_02581_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_267 ();
 sky130_fd_sc_hd__nand2_8 _09019_ (.A(_02595_),
    .B(_03367_),
    .Y(_03500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_266 ();
 sky130_fd_sc_hd__and3_1 _09021_ (.A(net191),
    .B(net97),
    .C(_03500_),
    .X(_03502_));
 sky130_fd_sc_hd__a21oi_1 _09022_ (.A1(_02588_),
    .A2(_03495_),
    .B1(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__o21ai_0 _09023_ (.A1(_02560_),
    .A2(_03496_),
    .B1(_03503_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _09024_ (.A(_02636_),
    .B(_03495_),
    .Y(_03504_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_265 ();
 sky130_fd_sc_hd__nand2_1 _09026_ (.A(net1267),
    .B(_03500_),
    .Y(_03506_));
 sky130_fd_sc_hd__a21oi_1 _09027_ (.A1(_03504_),
    .A2(_03506_),
    .B1(net108),
    .Y(_00673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_264 ();
 sky130_fd_sc_hd__nand2_1 _09029_ (.A(net1052),
    .B(_03500_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand2_1 _09030_ (.A(_02683_),
    .B(_03495_),
    .Y(_03509_));
 sky130_fd_sc_hd__a21oi_1 _09031_ (.A1(_03508_),
    .A2(_03509_),
    .B1(net109),
    .Y(_00674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_263 ();
 sky130_fd_sc_hd__nand3_1 _09033_ (.A(net1691),
    .B(net96),
    .C(_03500_),
    .Y(_03511_));
 sky130_fd_sc_hd__o21ai_0 _09034_ (.A1(_02713_),
    .A2(_03500_),
    .B1(_03511_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_02748_),
    .B(_03495_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(net1361),
    .B(_03500_),
    .Y(_03513_));
 sky130_fd_sc_hd__a21oi_1 _09037_ (.A1(_03512_),
    .A2(_03513_),
    .B1(net109),
    .Y(_00676_));
 sky130_fd_sc_hd__nand3_1 _09038_ (.A(net1419),
    .B(net97),
    .C(_03500_),
    .Y(_03514_));
 sky130_fd_sc_hd__o21ai_0 _09039_ (.A1(_02766_),
    .A2(_03500_),
    .B1(_03514_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand3_1 _09040_ (.A(net1371),
    .B(net97),
    .C(_03500_),
    .Y(_03515_));
 sky130_fd_sc_hd__o21ai_0 _09041_ (.A1(_02784_),
    .A2(_03500_),
    .B1(_03515_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand3_1 _09042_ (.A(net1398),
    .B(net97),
    .C(_03500_),
    .Y(_03516_));
 sky130_fd_sc_hd__o21ai_0 _09043_ (.A1(_02809_),
    .A2(_03500_),
    .B1(_03516_),
    .Y(_00679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_261 ();
 sky130_fd_sc_hd__nand3_1 _09046_ (.A(net1512),
    .B(net97),
    .C(_03500_),
    .Y(_03519_));
 sky130_fd_sc_hd__o221ai_1 _09047_ (.A1(_02834_),
    .A2(_03500_),
    .B1(_03496_),
    .B2(_02832_),
    .C1(_03519_),
    .Y(_00680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__and3_1 _09049_ (.A(net1759),
    .B(_02586_),
    .C(_03500_),
    .X(_03521_));
 sky130_fd_sc_hd__a31o_1 _09050_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03495_),
    .B1(_03521_),
    .X(_00681_));
 sky130_fd_sc_hd__and3_1 _09051_ (.A(net1811),
    .B(net97),
    .C(_03500_),
    .X(_03522_));
 sky130_fd_sc_hd__a21oi_1 _09052_ (.A1(_02884_),
    .A2(_03495_),
    .B1(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__o21ai_0 _09053_ (.A1(_02882_),
    .A2(_03496_),
    .B1(_03523_),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_1 _09054_ (.A(net171),
    .B(_03500_),
    .Y(_03524_));
 sky130_fd_sc_hd__o211ai_1 _09055_ (.A1(_02889_),
    .A2(_03500_),
    .B1(_03524_),
    .C1(_02586_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand3_1 _09056_ (.A(net1591),
    .B(net96),
    .C(_03500_),
    .Y(_03525_));
 sky130_fd_sc_hd__o221ai_1 _09057_ (.A1(_02909_),
    .A2(_03500_),
    .B1(_03496_),
    .B2(_02908_),
    .C1(_03525_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand3_1 _09058_ (.A(net1622),
    .B(_02586_),
    .C(_03500_),
    .Y(_03526_));
 sky130_fd_sc_hd__o221ai_1 _09059_ (.A1(_02936_),
    .A2(_03500_),
    .B1(_03496_),
    .B2(_02934_),
    .C1(_03526_),
    .Y(_00685_));
 sky130_fd_sc_hd__and3_1 _09060_ (.A(net1823),
    .B(_02586_),
    .C(_03500_),
    .X(_03527_));
 sky130_fd_sc_hd__a21oi_1 _09061_ (.A1(_02961_),
    .A2(_03495_),
    .B1(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21ai_0 _09062_ (.A1(_02959_),
    .A2(_03496_),
    .B1(_03528_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3_1 _09063_ (.A(net1665),
    .B(_02586_),
    .C(_03500_),
    .Y(_03529_));
 sky130_fd_sc_hd__o221ai_1 _09064_ (.A1(_02984_),
    .A2(_03500_),
    .B1(_03496_),
    .B2(_02983_),
    .C1(_03529_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _09065_ (.A(_03009_),
    .B(_03495_),
    .Y(_03530_));
 sky130_fd_sc_hd__nand2_1 _09066_ (.A(net1309),
    .B(_03500_),
    .Y(_03531_));
 sky130_fd_sc_hd__a21oi_1 _09067_ (.A1(_03530_),
    .A2(_03531_),
    .B1(net109),
    .Y(_00688_));
 sky130_fd_sc_hd__nor2_1 _09068_ (.A(_01035_),
    .B(_03500_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(_03031_),
    .B(_03495_),
    .Y(_03533_));
 sky130_fd_sc_hd__o21ai_0 _09070_ (.A1(net1704),
    .A2(_03495_),
    .B1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a311oi_1 _09071_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03532_),
    .B1(_03534_),
    .C1(net108),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _09072_ (.A(_03053_),
    .B(_03495_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(net1360),
    .B(_03500_),
    .Y(_03536_));
 sky130_fd_sc_hd__a21oi_1 _09074_ (.A1(_03535_),
    .A2(_03536_),
    .B1(net109),
    .Y(_00690_));
 sky130_fd_sc_hd__nand3_1 _09075_ (.A(net1597),
    .B(_02586_),
    .C(_03500_),
    .Y(_03537_));
 sky130_fd_sc_hd__o221ai_1 _09076_ (.A1(_03076_),
    .A2(_03500_),
    .B1(_03496_),
    .B2(_03074_),
    .C1(_03537_),
    .Y(_00691_));
 sky130_fd_sc_hd__and3_1 _09077_ (.A(net1824),
    .B(net97),
    .C(_03500_),
    .X(_03538_));
 sky130_fd_sc_hd__a21oi_1 _09078_ (.A1(_03100_),
    .A2(_03495_),
    .B1(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__o21ai_0 _09079_ (.A1(_03098_),
    .A2(_03496_),
    .B1(_03539_),
    .Y(_00692_));
 sky130_fd_sc_hd__a2111oi_0 _09080_ (.A1(net98),
    .A2(_03117_),
    .B1(_03500_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _09081_ (.A(net1559),
    .B(_03495_),
    .Y(_03541_));
 sky130_fd_sc_hd__a2111oi_0 _09082_ (.A1(_03104_),
    .A2(_03495_),
    .B1(_03540_),
    .C1(_03541_),
    .D1(net108),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _09083_ (.A(net168),
    .B(_03500_),
    .Y(_03542_));
 sky130_fd_sc_hd__o211ai_1 _09084_ (.A1(_03144_),
    .A2(_03500_),
    .B1(_03542_),
    .C1(_02586_),
    .Y(_00694_));
 sky130_fd_sc_hd__and3_1 _09085_ (.A(net1827),
    .B(_02586_),
    .C(_03500_),
    .X(_03543_));
 sky130_fd_sc_hd__a21oi_1 _09086_ (.A1(_03163_),
    .A2(_03495_),
    .B1(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__o21ai_0 _09087_ (.A1(_03161_),
    .A2(_03496_),
    .B1(_03544_),
    .Y(_00695_));
 sky130_fd_sc_hd__and3_1 _09088_ (.A(net1785),
    .B(net97),
    .C(_03500_),
    .X(_03545_));
 sky130_fd_sc_hd__a21oi_1 _09089_ (.A1(_03191_),
    .A2(_03495_),
    .B1(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__o21ai_0 _09090_ (.A1(_03189_),
    .A2(_03496_),
    .B1(_03546_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(net186),
    .B(_03500_),
    .Y(_03547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__o211ai_1 _09093_ (.A1(_03201_),
    .A2(_03500_),
    .B1(_03547_),
    .C1(net96),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_03210_),
    .B(_03495_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _09095_ (.A(net166),
    .B(_03500_),
    .Y(_03550_));
 sky130_fd_sc_hd__a21oi_1 _09096_ (.A1(_03549_),
    .A2(_03550_),
    .B1(net110),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _09097_ (.A(_03219_),
    .B(_03495_),
    .Y(_03551_));
 sky130_fd_sc_hd__nand2_1 _09098_ (.A(net180),
    .B(_03500_),
    .Y(_03552_));
 sky130_fd_sc_hd__a21oi_1 _09099_ (.A1(_03551_),
    .A2(_03552_),
    .B1(net110),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(_03227_),
    .B(_03495_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(net165),
    .B(_03500_),
    .Y(_03554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__a21oi_1 _09103_ (.A1(_03553_),
    .A2(_03554_),
    .B1(net110),
    .Y(_00700_));
 sky130_fd_sc_hd__nand3_1 _09104_ (.A(net504),
    .B(net96),
    .C(_03500_),
    .Y(_03556_));
 sky130_fd_sc_hd__o31ai_1 _09105_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03500_),
    .B1(_03556_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand3_1 _09106_ (.A(net195),
    .B(net96),
    .C(_03500_),
    .Y(_03557_));
 sky130_fd_sc_hd__o21ai_0 _09107_ (.A1(_03251_),
    .A2(_03500_),
    .B1(_03557_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand3_1 _09108_ (.A(net172),
    .B(net96),
    .C(_03500_),
    .Y(_03558_));
 sky130_fd_sc_hd__o31ai_1 _09109_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03500_),
    .B1(_03558_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_8 _09110_ (.A(_03269_),
    .B(_03367_),
    .Y(_03559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__a21oi_1 _09114_ (.A1(net1475),
    .A2(_03559_),
    .B1(CPU_reset_a3),
    .Y(_03563_));
 sky130_fd_sc_hd__o21ai_0 _09115_ (.A1(_03265_),
    .A2(_03559_),
    .B1(_03563_),
    .Y(_00704_));
 sky130_fd_sc_hd__nor2_8 _09116_ (.A(_03277_),
    .B(_03358_),
    .Y(_03564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 ();
 sky130_fd_sc_hd__nand2_1 _09118_ (.A(_02636_),
    .B(_03564_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_1 _09119_ (.A(net1278),
    .B(_03559_),
    .Y(_03567_));
 sky130_fd_sc_hd__a21oi_1 _09120_ (.A1(_03566_),
    .A2(_03567_),
    .B1(net108),
    .Y(_00705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 ();
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(net1335),
    .B(_03559_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _09123_ (.A(_02683_),
    .B(_03564_),
    .Y(_03570_));
 sky130_fd_sc_hd__a21oi_1 _09124_ (.A1(_03569_),
    .A2(_03570_),
    .B1(net109),
    .Y(_00706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__nand3_1 _09126_ (.A(net1564),
    .B(net96),
    .C(_03559_),
    .Y(_03572_));
 sky130_fd_sc_hd__o21ai_0 _09127_ (.A1(_02713_),
    .A2(_03559_),
    .B1(_03572_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_02748_),
    .B(_03564_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _09129_ (.A(net1235),
    .B(_03559_),
    .Y(_03574_));
 sky130_fd_sc_hd__a21oi_1 _09130_ (.A1(_03573_),
    .A2(_03574_),
    .B1(net109),
    .Y(_00708_));
 sky130_fd_sc_hd__nand3_1 _09131_ (.A(net1482),
    .B(net97),
    .C(_03559_),
    .Y(_03575_));
 sky130_fd_sc_hd__o21ai_0 _09132_ (.A1(_02766_),
    .A2(_03559_),
    .B1(_03575_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand3_1 _09133_ (.A(net1399),
    .B(net97),
    .C(_03559_),
    .Y(_03576_));
 sky130_fd_sc_hd__o21ai_0 _09134_ (.A1(_02784_),
    .A2(_03559_),
    .B1(_03576_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand3_1 _09135_ (.A(net1401),
    .B(net97),
    .C(_03559_),
    .Y(_03577_));
 sky130_fd_sc_hd__o21ai_0 _09136_ (.A1(_02809_),
    .A2(_03559_),
    .B1(_03577_),
    .Y(_00711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__nand2_8 _09138_ (.A(_02581_),
    .B(_03564_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand3_1 _09139_ (.A(net1498),
    .B(net97),
    .C(_03559_),
    .Y(_03580_));
 sky130_fd_sc_hd__o221ai_1 _09140_ (.A1(_02834_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_02832_),
    .C1(_03580_),
    .Y(_00712_));
 sky130_fd_sc_hd__and3_1 _09141_ (.A(net1767),
    .B(_02586_),
    .C(_03559_),
    .X(_03581_));
 sky130_fd_sc_hd__a31o_1 _09142_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03564_),
    .B1(_03581_),
    .X(_00713_));
 sky130_fd_sc_hd__and3_1 _09143_ (.A(net1773),
    .B(_02586_),
    .C(_03559_),
    .X(_03582_));
 sky130_fd_sc_hd__a21oi_1 _09144_ (.A1(_02884_),
    .A2(_03564_),
    .B1(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__o21ai_0 _09145_ (.A1(_02882_),
    .A2(_03579_),
    .B1(_03583_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _09146_ (.A(net1440),
    .B(_03559_),
    .Y(_03584_));
 sky130_fd_sc_hd__o211ai_1 _09147_ (.A1(_02889_),
    .A2(_03559_),
    .B1(_03584_),
    .C1(_02586_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand3_1 _09148_ (.A(net1653),
    .B(net97),
    .C(_03559_),
    .Y(_03585_));
 sky130_fd_sc_hd__o221ai_1 _09149_ (.A1(_02909_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_02908_),
    .C1(_03585_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand3_1 _09150_ (.A(net1636),
    .B(_02586_),
    .C(_03559_),
    .Y(_03586_));
 sky130_fd_sc_hd__o221ai_1 _09151_ (.A1(_02936_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_02934_),
    .C1(_03586_),
    .Y(_00717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__and3_1 _09153_ (.A(net1800),
    .B(_02586_),
    .C(_03559_),
    .X(_03588_));
 sky130_fd_sc_hd__a21oi_1 _09154_ (.A1(_02961_),
    .A2(_03564_),
    .B1(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__o21ai_0 _09155_ (.A1(_02959_),
    .A2(_03579_),
    .B1(_03589_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand3_1 _09156_ (.A(net1541),
    .B(_02586_),
    .C(_03559_),
    .Y(_03590_));
 sky130_fd_sc_hd__o221ai_1 _09157_ (.A1(_02984_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_02983_),
    .C1(_03590_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_03009_),
    .B(_03564_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand2_1 _09159_ (.A(net1326),
    .B(_03559_),
    .Y(_03592_));
 sky130_fd_sc_hd__a21oi_1 _09160_ (.A1(_03591_),
    .A2(_03592_),
    .B1(net109),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_1 _09161_ (.A(_01035_),
    .B(_03559_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _09162_ (.A(_03031_),
    .B(_03564_),
    .Y(_03594_));
 sky130_fd_sc_hd__o21ai_0 _09163_ (.A1(net1696),
    .A2(_03564_),
    .B1(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__a311oi_1 _09164_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03593_),
    .B1(_03595_),
    .C1(net108),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_1 _09165_ (.A(_03053_),
    .B(_03564_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _09166_ (.A(net1336),
    .B(_03559_),
    .Y(_03597_));
 sky130_fd_sc_hd__a21oi_1 _09167_ (.A1(_03596_),
    .A2(_03597_),
    .B1(net109),
    .Y(_00722_));
 sky130_fd_sc_hd__nand3_1 _09168_ (.A(net1522),
    .B(_02586_),
    .C(_03559_),
    .Y(_03598_));
 sky130_fd_sc_hd__o221ai_1 _09169_ (.A1(_03076_),
    .A2(_03559_),
    .B1(_03579_),
    .B2(_03074_),
    .C1(_03598_),
    .Y(_00723_));
 sky130_fd_sc_hd__and3_1 _09170_ (.A(net1784),
    .B(_02586_),
    .C(_03559_),
    .X(_03599_));
 sky130_fd_sc_hd__a21oi_1 _09171_ (.A1(_03100_),
    .A2(_03564_),
    .B1(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__o21ai_0 _09172_ (.A1(_03098_),
    .A2(_03579_),
    .B1(_03600_),
    .Y(_00724_));
 sky130_fd_sc_hd__a2111oi_0 _09173_ (.A1(net98),
    .A2(_03117_),
    .B1(_03559_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03601_));
 sky130_fd_sc_hd__nor2_1 _09174_ (.A(net1593),
    .B(_03564_),
    .Y(_03602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_249 ();
 sky130_fd_sc_hd__a2111oi_0 _09176_ (.A1(_03104_),
    .A2(_03564_),
    .B1(_03601_),
    .C1(_03602_),
    .D1(net108),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_1 _09177_ (.A(net1552),
    .B(_03559_),
    .Y(_03604_));
 sky130_fd_sc_hd__o211ai_1 _09178_ (.A1(_03144_),
    .A2(_03559_),
    .B1(_03604_),
    .C1(net96),
    .Y(_00726_));
 sky130_fd_sc_hd__and3_1 _09179_ (.A(net1834),
    .B(_02586_),
    .C(_03559_),
    .X(_03605_));
 sky130_fd_sc_hd__a21oi_1 _09180_ (.A1(_03163_),
    .A2(_03564_),
    .B1(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__o21ai_0 _09181_ (.A1(_03161_),
    .A2(_03579_),
    .B1(_03606_),
    .Y(_00727_));
 sky130_fd_sc_hd__and3_1 _09182_ (.A(net1752),
    .B(net97),
    .C(_03559_),
    .X(_03607_));
 sky130_fd_sc_hd__a21oi_1 _09183_ (.A1(_03191_),
    .A2(_03564_),
    .B1(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21ai_0 _09184_ (.A1(_03189_),
    .A2(_03579_),
    .B1(_03608_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _09185_ (.A(net1438),
    .B(_03559_),
    .Y(_03609_));
 sky130_fd_sc_hd__o211ai_1 _09186_ (.A1(_03201_),
    .A2(_03559_),
    .B1(_03609_),
    .C1(net96),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(_03210_),
    .B(_03564_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand2_1 _09188_ (.A(net1271),
    .B(_03559_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21oi_1 _09189_ (.A1(_03610_),
    .A2(_03611_),
    .B1(net110),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_03219_),
    .B(_03564_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _09191_ (.A(net1275),
    .B(_03559_),
    .Y(_03613_));
 sky130_fd_sc_hd__a21oi_1 _09192_ (.A1(_03612_),
    .A2(_03613_),
    .B1(CPU_reset_a3),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _09193_ (.A(_03227_),
    .B(_03564_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(net1294),
    .B(_03559_),
    .Y(_03615_));
 sky130_fd_sc_hd__a21oi_1 _09195_ (.A1(_03614_),
    .A2(_03615_),
    .B1(net110),
    .Y(_00732_));
 sky130_fd_sc_hd__nand3_1 _09196_ (.A(net1468),
    .B(net96),
    .C(_03559_),
    .Y(_03616_));
 sky130_fd_sc_hd__o31ai_1 _09197_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03559_),
    .B1(_03616_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand3_1 _09198_ (.A(net1355),
    .B(net96),
    .C(_03559_),
    .Y(_03617_));
 sky130_fd_sc_hd__o21ai_0 _09199_ (.A1(_03251_),
    .A2(_03559_),
    .B1(_03617_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand3_1 _09200_ (.A(net1412),
    .B(net96),
    .C(_03559_),
    .Y(_03618_));
 sky130_fd_sc_hd__o31ai_1 _09201_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03559_),
    .B1(_03618_),
    .Y(_00735_));
 sky130_fd_sc_hd__nor3_1 _09202_ (.A(\CPU_rd_a5[2] ),
    .B(\CPU_rd_a5[3] ),
    .C(_01036_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21oi_4 _09203_ (.A1(_01036_),
    .A2(_02571_),
    .B1(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_8 _09204_ (.A(_02593_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_8 _09205_ (.A(_03437_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_246 ();
 sky130_fd_sc_hd__a21oi_1 _09209_ (.A1(net1485),
    .A2(_03622_),
    .B1(net108),
    .Y(_03626_));
 sky130_fd_sc_hd__o21ai_0 _09210_ (.A1(_03265_),
    .A2(_03622_),
    .B1(_03626_),
    .Y(_00736_));
 sky130_fd_sc_hd__nor3_4 _09211_ (.A(_02593_),
    .B(_03430_),
    .C(_03620_),
    .Y(_03627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_245 ();
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(_02636_),
    .B(_03627_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand2_1 _09214_ (.A(net1287),
    .B(_03622_),
    .Y(_03630_));
 sky130_fd_sc_hd__a21oi_1 _09215_ (.A1(_03629_),
    .A2(_03630_),
    .B1(net108),
    .Y(_00737_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_244 ();
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(net1190),
    .B(_03622_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_02683_),
    .B(net13),
    .Y(_03633_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_243 ();
 sky130_fd_sc_hd__a21oi_1 _09220_ (.A1(_03632_),
    .A2(_03633_),
    .B1(net109),
    .Y(_00738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_242 ();
 sky130_fd_sc_hd__nand3_1 _09222_ (.A(net1494),
    .B(net96),
    .C(_03622_),
    .Y(_03636_));
 sky130_fd_sc_hd__o21ai_0 _09223_ (.A1(_02713_),
    .A2(_03622_),
    .B1(_03636_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(_02748_),
    .B(net13),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2_1 _09225_ (.A(net1135),
    .B(_03622_),
    .Y(_03638_));
 sky130_fd_sc_hd__a21oi_1 _09226_ (.A1(_03637_),
    .A2(_03638_),
    .B1(net109),
    .Y(_00740_));
 sky130_fd_sc_hd__nand3_1 _09227_ (.A(net1467),
    .B(net97),
    .C(_03622_),
    .Y(_03639_));
 sky130_fd_sc_hd__o21ai_0 _09228_ (.A1(_02766_),
    .A2(_03622_),
    .B1(_03639_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand3_1 _09229_ (.A(net1670),
    .B(net97),
    .C(_03622_),
    .Y(_03640_));
 sky130_fd_sc_hd__o21ai_0 _09230_ (.A1(_02784_),
    .A2(_03622_),
    .B1(_03640_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand3_1 _09231_ (.A(net1442),
    .B(net97),
    .C(_03622_),
    .Y(_03641_));
 sky130_fd_sc_hd__o21ai_0 _09232_ (.A1(_02809_),
    .A2(_03622_),
    .B1(_03641_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_8 _09233_ (.A(_02581_),
    .B(net13),
    .Y(_03642_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_241 ();
 sky130_fd_sc_hd__nand3_1 _09235_ (.A(net1644),
    .B(net97),
    .C(_03622_),
    .Y(_03644_));
 sky130_fd_sc_hd__o221ai_1 _09236_ (.A1(_02834_),
    .A2(_03622_),
    .B1(_03642_),
    .B2(_02832_),
    .C1(_03644_),
    .Y(_00744_));
 sky130_fd_sc_hd__and3_1 _09237_ (.A(net1795),
    .B(_02586_),
    .C(_03622_),
    .X(_03645_));
 sky130_fd_sc_hd__a31o_1 _09238_ (.A1(_02854_),
    .A2(_02856_),
    .A3(net13),
    .B1(_03645_),
    .X(_00745_));
 sky130_fd_sc_hd__and3_1 _09239_ (.A(net1837),
    .B(net97),
    .C(_03622_),
    .X(_03646_));
 sky130_fd_sc_hd__a21oi_1 _09240_ (.A1(_02884_),
    .A2(_03627_),
    .B1(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__o21ai_0 _09241_ (.A1(_02882_),
    .A2(_03642_),
    .B1(_03647_),
    .Y(_00746_));
 sky130_fd_sc_hd__nor2_1 _09242_ (.A(_02889_),
    .B(_03622_),
    .Y(_03648_));
 sky130_fd_sc_hd__a21oi_1 _09243_ (.A1(net1632),
    .A2(_03622_),
    .B1(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__nor2_1 _09244_ (.A(CPU_reset_a3),
    .B(_03649_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand3_1 _09245_ (.A(net1586),
    .B(net97),
    .C(_03622_),
    .Y(_03650_));
 sky130_fd_sc_hd__o221ai_1 _09246_ (.A1(_02909_),
    .A2(_03622_),
    .B1(_03642_),
    .B2(_02908_),
    .C1(_03650_),
    .Y(_00748_));
 sky130_fd_sc_hd__nand3_1 _09247_ (.A(net1682),
    .B(net97),
    .C(_03622_),
    .Y(_03651_));
 sky130_fd_sc_hd__o221ai_1 _09248_ (.A1(_02936_),
    .A2(_03622_),
    .B1(_03642_),
    .B2(_02934_),
    .C1(_03651_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand3_1 _09249_ (.A(net1471),
    .B(_02586_),
    .C(_03622_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(_02961_),
    .B(net13),
    .Y(_03653_));
 sky130_fd_sc_hd__o211ai_1 _09251_ (.A1(_02959_),
    .A2(_03642_),
    .B1(_03652_),
    .C1(_03653_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand3_1 _09252_ (.A(net1640),
    .B(net97),
    .C(_03622_),
    .Y(_03654_));
 sky130_fd_sc_hd__o221ai_1 _09253_ (.A1(_02984_),
    .A2(_03622_),
    .B1(_03642_),
    .B2(_02983_),
    .C1(_03654_),
    .Y(_00751_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(_03009_),
    .B(net13),
    .Y(_03655_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(net1242),
    .B(_03622_),
    .Y(_03656_));
 sky130_fd_sc_hd__a21oi_1 _09256_ (.A1(_03655_),
    .A2(_03656_),
    .B1(net109),
    .Y(_00752_));
 sky130_fd_sc_hd__nor2_1 _09257_ (.A(_01035_),
    .B(_03622_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand2_1 _09258_ (.A(_03031_),
    .B(_03627_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_0 _09259_ (.A1(net1695),
    .A2(_03627_),
    .B1(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__a311oi_1 _09260_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03657_),
    .B1(_03659_),
    .C1(net108),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_03053_),
    .B(net13),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(net1333),
    .B(_03622_),
    .Y(_03661_));
 sky130_fd_sc_hd__a21oi_1 _09263_ (.A1(_03660_),
    .A2(_03661_),
    .B1(net109),
    .Y(_00754_));
 sky130_fd_sc_hd__nand3_1 _09264_ (.A(net1625),
    .B(_02586_),
    .C(_03622_),
    .Y(_03662_));
 sky130_fd_sc_hd__o221ai_1 _09265_ (.A1(_03076_),
    .A2(_03622_),
    .B1(_03642_),
    .B2(_03074_),
    .C1(_03662_),
    .Y(_00755_));
 sky130_fd_sc_hd__and3_1 _09266_ (.A(net1829),
    .B(_02586_),
    .C(_03622_),
    .X(_03663_));
 sky130_fd_sc_hd__a21oi_1 _09267_ (.A1(_03100_),
    .A2(net13),
    .B1(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__o21ai_0 _09268_ (.A1(_03098_),
    .A2(_03642_),
    .B1(_03664_),
    .Y(_00756_));
 sky130_fd_sc_hd__a2111oi_0 _09269_ (.A1(net98),
    .A2(_03117_),
    .B1(_03622_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03665_));
 sky130_fd_sc_hd__nor2_1 _09270_ (.A(net1633),
    .B(_03627_),
    .Y(_03666_));
 sky130_fd_sc_hd__a2111oi_0 _09271_ (.A1(_03104_),
    .A2(_03627_),
    .B1(_03665_),
    .C1(_03666_),
    .D1(net108),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _09272_ (.A(_03144_),
    .B(_03622_),
    .Y(_03667_));
 sky130_fd_sc_hd__a21oi_1 _09273_ (.A1(net1579),
    .A2(_03622_),
    .B1(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__nor2_1 _09274_ (.A(net110),
    .B(_03668_),
    .Y(_00758_));
 sky130_fd_sc_hd__and3_1 _09275_ (.A(net1816),
    .B(_02586_),
    .C(_03622_),
    .X(_03669_));
 sky130_fd_sc_hd__a21oi_1 _09276_ (.A1(_03163_),
    .A2(net13),
    .B1(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__o21ai_0 _09277_ (.A1(_03161_),
    .A2(_03642_),
    .B1(_03670_),
    .Y(_00759_));
 sky130_fd_sc_hd__and3_1 _09278_ (.A(net1809),
    .B(net97),
    .C(_03622_),
    .X(_03671_));
 sky130_fd_sc_hd__a21oi_1 _09279_ (.A1(_03191_),
    .A2(net13),
    .B1(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__o21ai_0 _09280_ (.A1(_03189_),
    .A2(_03642_),
    .B1(_03672_),
    .Y(_00760_));
 sky130_fd_sc_hd__nor2_1 _09281_ (.A(_03201_),
    .B(_03622_),
    .Y(_03673_));
 sky130_fd_sc_hd__a21oi_1 _09282_ (.A1(net1599),
    .A2(_03622_),
    .B1(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__nor2_1 _09283_ (.A(CPU_reset_a3),
    .B(_03674_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _09284_ (.A(_03210_),
    .B(_03627_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _09285_ (.A(net1280),
    .B(_03622_),
    .Y(_03676_));
 sky130_fd_sc_hd__a21oi_1 _09286_ (.A1(_03675_),
    .A2(_03676_),
    .B1(net110),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_03219_),
    .B(_03627_),
    .Y(_03677_));
 sky130_fd_sc_hd__nand2_1 _09288_ (.A(net1138),
    .B(_03622_),
    .Y(_03678_));
 sky130_fd_sc_hd__a21oi_1 _09289_ (.A1(_03677_),
    .A2(_03678_),
    .B1(CPU_reset_a3),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(_03227_),
    .B(net13),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(net1289),
    .B(_03622_),
    .Y(_03680_));
 sky130_fd_sc_hd__a21oi_1 _09292_ (.A1(_03679_),
    .A2(_03680_),
    .B1(net110),
    .Y(_00764_));
 sky130_fd_sc_hd__nand3_1 _09293_ (.A(net1472),
    .B(net96),
    .C(_03622_),
    .Y(_03681_));
 sky130_fd_sc_hd__o31ai_1 _09294_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03622_),
    .B1(_03681_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand3_1 _09295_ (.A(net1497),
    .B(net96),
    .C(_03622_),
    .Y(_03682_));
 sky130_fd_sc_hd__o21ai_0 _09296_ (.A1(_03251_),
    .A2(_03622_),
    .B1(_03682_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand3_1 _09297_ (.A(net1396),
    .B(net96),
    .C(_03622_),
    .Y(_03683_));
 sky130_fd_sc_hd__o31ai_1 _09298_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03622_),
    .B1(_03683_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor3_4 _09299_ (.A(_02593_),
    .B(_02594_),
    .C(_03620_),
    .Y(_03684_));
 sky130_fd_sc_hd__nand2_8 _09300_ (.A(_02581_),
    .B(net12),
    .Y(_03685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_238 ();
 sky130_fd_sc_hd__nand2_8 _09304_ (.A(_02578_),
    .B(_03621_),
    .Y(_03689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_237 ();
 sky130_fd_sc_hd__and3_1 _09306_ (.A(net1826),
    .B(net96),
    .C(_03689_),
    .X(_03691_));
 sky130_fd_sc_hd__a21oi_1 _09307_ (.A1(_02588_),
    .A2(net12),
    .B1(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__o21ai_0 _09308_ (.A1(_02560_),
    .A2(_03685_),
    .B1(_03692_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_02636_),
    .B(_03684_),
    .Y(_03693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_236 ();
 sky130_fd_sc_hd__nand2_1 _09311_ (.A(net1297),
    .B(_03689_),
    .Y(_03695_));
 sky130_fd_sc_hd__a21oi_1 _09312_ (.A1(_03693_),
    .A2(_03695_),
    .B1(net108),
    .Y(_00769_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_235 ();
 sky130_fd_sc_hd__nand2_1 _09314_ (.A(net1173),
    .B(_03689_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_1 _09315_ (.A(_02683_),
    .B(net12),
    .Y(_03698_));
 sky130_fd_sc_hd__a21oi_1 _09316_ (.A1(_03697_),
    .A2(_03698_),
    .B1(net109),
    .Y(_00770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_232 ();
 sky130_fd_sc_hd__nand3_1 _09320_ (.A(net1635),
    .B(net96),
    .C(_03689_),
    .Y(_03702_));
 sky130_fd_sc_hd__o21ai_0 _09321_ (.A1(_02713_),
    .A2(_03689_),
    .B1(_03702_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _09322_ (.A(net1113),
    .B(_03689_),
    .Y(_03703_));
 sky130_fd_sc_hd__nand2_1 _09323_ (.A(_02748_),
    .B(net12),
    .Y(_03704_));
 sky130_fd_sc_hd__a21oi_1 _09324_ (.A1(_03703_),
    .A2(_03704_),
    .B1(net109),
    .Y(_00772_));
 sky130_fd_sc_hd__nand3_1 _09325_ (.A(net1397),
    .B(net97),
    .C(_03689_),
    .Y(_03705_));
 sky130_fd_sc_hd__o21ai_0 _09326_ (.A1(_02766_),
    .A2(_03689_),
    .B1(_03705_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand3_1 _09327_ (.A(net1568),
    .B(net97),
    .C(_03689_),
    .Y(_03706_));
 sky130_fd_sc_hd__o21ai_0 _09328_ (.A1(_02784_),
    .A2(_03689_),
    .B1(_03706_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand3_1 _09329_ (.A(net1439),
    .B(net97),
    .C(_03689_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ai_0 _09330_ (.A1(_02809_),
    .A2(_03689_),
    .B1(_03707_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand3_1 _09331_ (.A(net1641),
    .B(net97),
    .C(_03689_),
    .Y(_03708_));
 sky130_fd_sc_hd__o221ai_1 _09332_ (.A1(_02834_),
    .A2(_03689_),
    .B1(_03685_),
    .B2(_02832_),
    .C1(_03708_),
    .Y(_00776_));
 sky130_fd_sc_hd__and3_1 _09333_ (.A(net1770),
    .B(_02586_),
    .C(_03689_),
    .X(_03709_));
 sky130_fd_sc_hd__a31o_1 _09334_ (.A1(_02854_),
    .A2(_02856_),
    .A3(net12),
    .B1(_03709_),
    .X(_00777_));
 sky130_fd_sc_hd__and3_1 _09335_ (.A(net1796),
    .B(net97),
    .C(_03689_),
    .X(_03710_));
 sky130_fd_sc_hd__a21oi_1 _09336_ (.A1(_02884_),
    .A2(net12),
    .B1(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__o21ai_0 _09337_ (.A1(_02882_),
    .A2(_03685_),
    .B1(_03711_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _09338_ (.A(net1477),
    .B(_03689_),
    .Y(_03712_));
 sky130_fd_sc_hd__o211ai_1 _09339_ (.A1(_02889_),
    .A2(_03689_),
    .B1(_03712_),
    .C1(_02586_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand3_1 _09340_ (.A(net1575),
    .B(net96),
    .C(_03689_),
    .Y(_03713_));
 sky130_fd_sc_hd__o221ai_1 _09341_ (.A1(_02909_),
    .A2(_03689_),
    .B1(_03685_),
    .B2(_02908_),
    .C1(_03713_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand3_1 _09342_ (.A(net1539),
    .B(net96),
    .C(_03689_),
    .Y(_03714_));
 sky130_fd_sc_hd__o221ai_1 _09343_ (.A1(_02936_),
    .A2(_03689_),
    .B1(_03685_),
    .B2(_02934_),
    .C1(_03714_),
    .Y(_00781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_231 ();
 sky130_fd_sc_hd__and3_1 _09345_ (.A(net1813),
    .B(_02586_),
    .C(_03689_),
    .X(_03716_));
 sky130_fd_sc_hd__a21oi_1 _09346_ (.A1(_02961_),
    .A2(net12),
    .B1(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__o21ai_0 _09347_ (.A1(_02959_),
    .A2(_03685_),
    .B1(_03717_),
    .Y(_00782_));
 sky130_fd_sc_hd__nand3_1 _09348_ (.A(net1555),
    .B(net97),
    .C(_03689_),
    .Y(_03718_));
 sky130_fd_sc_hd__o221ai_1 _09349_ (.A1(_02984_),
    .A2(_03689_),
    .B1(_03685_),
    .B2(_02983_),
    .C1(_03718_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand2_1 _09350_ (.A(net1215),
    .B(_03689_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(_03009_),
    .B(net12),
    .Y(_03720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_230 ();
 sky130_fd_sc_hd__a21oi_1 _09353_ (.A1(_03719_),
    .A2(_03720_),
    .B1(net109),
    .Y(_00784_));
 sky130_fd_sc_hd__nor2_1 _09354_ (.A(_01035_),
    .B(_03689_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _09355_ (.A(_03031_),
    .B(_03684_),
    .Y(_03723_));
 sky130_fd_sc_hd__o21ai_0 _09356_ (.A1(net1702),
    .A2(_03684_),
    .B1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__a311oi_1 _09357_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03722_),
    .B1(_03724_),
    .C1(net108),
    .Y(_00785_));
 sky130_fd_sc_hd__nand2_1 _09358_ (.A(net1223),
    .B(_03689_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _09359_ (.A(_03053_),
    .B(net12),
    .Y(_03726_));
 sky130_fd_sc_hd__a21oi_1 _09360_ (.A1(_03725_),
    .A2(_03726_),
    .B1(net109),
    .Y(_00786_));
 sky130_fd_sc_hd__nand3_1 _09361_ (.A(net1687),
    .B(_02586_),
    .C(_03689_),
    .Y(_03727_));
 sky130_fd_sc_hd__o221ai_1 _09362_ (.A1(_03076_),
    .A2(_03689_),
    .B1(_03685_),
    .B2(_03074_),
    .C1(_03727_),
    .Y(_00787_));
 sky130_fd_sc_hd__and3_1 _09363_ (.A(net1844),
    .B(net97),
    .C(_03689_),
    .X(_03728_));
 sky130_fd_sc_hd__a21oi_1 _09364_ (.A1(_03100_),
    .A2(net12),
    .B1(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__o21ai_0 _09365_ (.A1(_03098_),
    .A2(_03685_),
    .B1(_03729_),
    .Y(_00788_));
 sky130_fd_sc_hd__a2111oi_0 _09366_ (.A1(net98),
    .A2(_03117_),
    .B1(_03689_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _09367_ (.A(net1611),
    .B(_03684_),
    .Y(_03731_));
 sky130_fd_sc_hd__a2111oi_0 _09368_ (.A1(_03104_),
    .A2(_03684_),
    .B1(_03730_),
    .C1(_03731_),
    .D1(net108),
    .Y(_00789_));
 sky130_fd_sc_hd__nor2_1 _09369_ (.A(_03144_),
    .B(_03689_),
    .Y(_03732_));
 sky130_fd_sc_hd__a21oi_1 _09370_ (.A1(net1561),
    .A2(_03689_),
    .B1(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _09371_ (.A(CPU_reset_a3),
    .B(_03733_),
    .Y(_00790_));
 sky130_fd_sc_hd__and3_1 _09372_ (.A(net1817),
    .B(_02586_),
    .C(_03689_),
    .X(_03734_));
 sky130_fd_sc_hd__a21oi_1 _09373_ (.A1(_03163_),
    .A2(net12),
    .B1(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__o21ai_0 _09374_ (.A1(_03161_),
    .A2(_03685_),
    .B1(_03735_),
    .Y(_00791_));
 sky130_fd_sc_hd__and3_1 _09375_ (.A(net1825),
    .B(net97),
    .C(_03689_),
    .X(_03736_));
 sky130_fd_sc_hd__a21oi_1 _09376_ (.A1(_03191_),
    .A2(net12),
    .B1(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__o21ai_0 _09377_ (.A1(_03189_),
    .A2(_03685_),
    .B1(_03737_),
    .Y(_00792_));
 sky130_fd_sc_hd__nor2_1 _09378_ (.A(_03201_),
    .B(_03689_),
    .Y(_03738_));
 sky130_fd_sc_hd__a21oi_1 _09379_ (.A1(net1667),
    .A2(_03689_),
    .B1(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _09380_ (.A(CPU_reset_a3),
    .B(_03739_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_03210_),
    .B(net12),
    .Y(_03740_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(net1276),
    .B(_03689_),
    .Y(_03741_));
 sky130_fd_sc_hd__a21oi_1 _09383_ (.A1(_03740_),
    .A2(_03741_),
    .B1(net110),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_03219_),
    .B(_03684_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(net1304),
    .B(_03689_),
    .Y(_03743_));
 sky130_fd_sc_hd__a21oi_1 _09386_ (.A1(_03742_),
    .A2(_03743_),
    .B1(CPU_reset_a3),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _09387_ (.A(_03227_),
    .B(net12),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(net1305),
    .B(_03689_),
    .Y(_03745_));
 sky130_fd_sc_hd__a21oi_1 _09389_ (.A1(_03744_),
    .A2(_03745_),
    .B1(net110),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_1 _09390_ (.A(net1479),
    .B(net96),
    .C(_03689_),
    .Y(_03746_));
 sky130_fd_sc_hd__o31ai_1 _09391_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03689_),
    .B1(_03746_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand3_1 _09392_ (.A(net1462),
    .B(net96),
    .C(_03689_),
    .Y(_03747_));
 sky130_fd_sc_hd__o21ai_0 _09393_ (.A1(_03251_),
    .A2(_03689_),
    .B1(_03747_),
    .Y(_00798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_229 ();
 sky130_fd_sc_hd__nand3_1 _09395_ (.A(net1466),
    .B(net96),
    .C(_03689_),
    .Y(_03749_));
 sky130_fd_sc_hd__o31ai_1 _09396_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03689_),
    .B1(_03749_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_8 _09397_ (.A(_03268_),
    .B(_03621_),
    .Y(_03750_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_226 ();
 sky130_fd_sc_hd__a21oi_1 _09401_ (.A1(net1483),
    .A2(_03750_),
    .B1(net108),
    .Y(_03754_));
 sky130_fd_sc_hd__o21ai_0 _09402_ (.A1(_03265_),
    .A2(_03750_),
    .B1(_03754_),
    .Y(_00800_));
 sky130_fd_sc_hd__and2_4 _09403_ (.A(_03268_),
    .B(_03621_),
    .X(_03755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_224 ();
 sky130_fd_sc_hd__nand2_1 _09406_ (.A(_02636_),
    .B(_03755_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _09407_ (.A(net1308),
    .B(_03750_),
    .Y(_03759_));
 sky130_fd_sc_hd__a21oi_1 _09408_ (.A1(_03758_),
    .A2(_03759_),
    .B1(net108),
    .Y(_00801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_223 ();
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(net1118),
    .B(_03750_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_1 _09411_ (.A(_02683_),
    .B(_03755_),
    .Y(_03762_));
 sky130_fd_sc_hd__a21oi_1 _09412_ (.A1(_03761_),
    .A2(_03762_),
    .B1(net109),
    .Y(_00802_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_222 ();
 sky130_fd_sc_hd__nand3_1 _09414_ (.A(net1441),
    .B(net96),
    .C(_03750_),
    .Y(_03764_));
 sky130_fd_sc_hd__o21ai_0 _09415_ (.A1(_02713_),
    .A2(_03750_),
    .B1(_03764_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_1 _09416_ (.A(_02748_),
    .B(_03755_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _09417_ (.A(net1186),
    .B(_03750_),
    .Y(_03766_));
 sky130_fd_sc_hd__a21oi_1 _09418_ (.A1(_03765_),
    .A2(_03766_),
    .B1(net109),
    .Y(_00804_));
 sky130_fd_sc_hd__nand3_1 _09419_ (.A(net1376),
    .B(net97),
    .C(_03750_),
    .Y(_03767_));
 sky130_fd_sc_hd__o21ai_0 _09420_ (.A1(_02766_),
    .A2(_03750_),
    .B1(_03767_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand3_1 _09421_ (.A(net1707),
    .B(net97),
    .C(_03750_),
    .Y(_03768_));
 sky130_fd_sc_hd__o21ai_0 _09422_ (.A1(_02784_),
    .A2(_03750_),
    .B1(_03768_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand3_1 _09423_ (.A(net1384),
    .B(net97),
    .C(_03750_),
    .Y(_03769_));
 sky130_fd_sc_hd__o21ai_0 _09424_ (.A1(_02809_),
    .A2(_03750_),
    .B1(_03769_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_8 _09425_ (.A(_02581_),
    .B(_03755_),
    .Y(_03770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_221 ();
 sky130_fd_sc_hd__nand3_1 _09427_ (.A(net1549),
    .B(net97),
    .C(_03750_),
    .Y(_03772_));
 sky130_fd_sc_hd__o221ai_1 _09428_ (.A1(_02834_),
    .A2(_03750_),
    .B1(_03770_),
    .B2(_02832_),
    .C1(_03772_),
    .Y(_00808_));
 sky130_fd_sc_hd__and3_1 _09429_ (.A(net1728),
    .B(_02586_),
    .C(_03750_),
    .X(_03773_));
 sky130_fd_sc_hd__a31o_1 _09430_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03755_),
    .B1(_03773_),
    .X(_00809_));
 sky130_fd_sc_hd__and3_1 _09431_ (.A(net1747),
    .B(net97),
    .C(_03750_),
    .X(_03774_));
 sky130_fd_sc_hd__a21oi_1 _09432_ (.A1(_02884_),
    .A2(_03755_),
    .B1(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__o21ai_0 _09433_ (.A1(_02882_),
    .A2(_03770_),
    .B1(_03775_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _09434_ (.A(net1490),
    .B(_03750_),
    .Y(_03776_));
 sky130_fd_sc_hd__o211ai_1 _09435_ (.A1(_02889_),
    .A2(_03750_),
    .B1(_03776_),
    .C1(_02586_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand3_1 _09436_ (.A(net1681),
    .B(net97),
    .C(_03750_),
    .Y(_03777_));
 sky130_fd_sc_hd__o221ai_1 _09437_ (.A1(_02909_),
    .A2(_03750_),
    .B1(_03770_),
    .B2(_02908_),
    .C1(_03777_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand3_1 _09438_ (.A(net1677),
    .B(_02586_),
    .C(_03750_),
    .Y(_03778_));
 sky130_fd_sc_hd__o221ai_1 _09439_ (.A1(_02936_),
    .A2(_03750_),
    .B1(_03770_),
    .B2(_02934_),
    .C1(_03778_),
    .Y(_00813_));
 sky130_fd_sc_hd__and3_1 _09440_ (.A(net1763),
    .B(_02586_),
    .C(_03750_),
    .X(_03779_));
 sky130_fd_sc_hd__a21oi_1 _09441_ (.A1(_02961_),
    .A2(_03755_),
    .B1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o21ai_0 _09442_ (.A1(_02959_),
    .A2(_03770_),
    .B1(_03780_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand3_1 _09443_ (.A(net1688),
    .B(_02586_),
    .C(_03750_),
    .Y(_03781_));
 sky130_fd_sc_hd__o221ai_1 _09444_ (.A1(_02984_),
    .A2(_03750_),
    .B1(_03770_),
    .B2(_02983_),
    .C1(_03781_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _09445_ (.A(_03009_),
    .B(_03755_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(net1170),
    .B(_03750_),
    .Y(_03783_));
 sky130_fd_sc_hd__a21oi_1 _09447_ (.A1(_03782_),
    .A2(_03783_),
    .B1(net109),
    .Y(_00816_));
 sky130_fd_sc_hd__nor2_1 _09448_ (.A(_01035_),
    .B(_03750_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _09449_ (.A(_03031_),
    .B(_03755_),
    .Y(_03785_));
 sky130_fd_sc_hd__o21ai_0 _09450_ (.A1(net1703),
    .A2(_03755_),
    .B1(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__a311oi_1 _09451_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03784_),
    .B1(_03786_),
    .C1(net108),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_03053_),
    .B(_03755_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(net1226),
    .B(_03750_),
    .Y(_03788_));
 sky130_fd_sc_hd__a21oi_1 _09454_ (.A1(_03787_),
    .A2(_03788_),
    .B1(net109),
    .Y(_00818_));
 sky130_fd_sc_hd__nand3_1 _09455_ (.A(net1639),
    .B(_02586_),
    .C(_03750_),
    .Y(_03789_));
 sky130_fd_sc_hd__o221ai_1 _09456_ (.A1(_03076_),
    .A2(_03750_),
    .B1(_03770_),
    .B2(_03074_),
    .C1(_03789_),
    .Y(_00819_));
 sky130_fd_sc_hd__and3_1 _09457_ (.A(net1775),
    .B(net97),
    .C(_03750_),
    .X(_03790_));
 sky130_fd_sc_hd__a21oi_1 _09458_ (.A1(_03100_),
    .A2(_03755_),
    .B1(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__o21ai_0 _09459_ (.A1(_03098_),
    .A2(_03770_),
    .B1(_03791_),
    .Y(_00820_));
 sky130_fd_sc_hd__a2111oi_0 _09460_ (.A1(net98),
    .A2(_03117_),
    .B1(_03750_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _09461_ (.A(net1637),
    .B(_03755_),
    .Y(_03793_));
 sky130_fd_sc_hd__a2111oi_0 _09462_ (.A1(_03104_),
    .A2(_03755_),
    .B1(_03792_),
    .C1(_03793_),
    .D1(net108),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_1 _09463_ (.A(_03144_),
    .B(_03750_),
    .Y(_03794_));
 sky130_fd_sc_hd__a21oi_1 _09464_ (.A1(net1627),
    .A2(_03750_),
    .B1(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(net110),
    .B(_03795_),
    .Y(_00822_));
 sky130_fd_sc_hd__and3_1 _09466_ (.A(net1749),
    .B(_02586_),
    .C(_03750_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_1 _09467_ (.A1(_03163_),
    .A2(_03755_),
    .B1(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__o21ai_0 _09468_ (.A1(_03161_),
    .A2(_03770_),
    .B1(_03797_),
    .Y(_00823_));
 sky130_fd_sc_hd__and3_1 _09469_ (.A(net1803),
    .B(net97),
    .C(_03750_),
    .X(_03798_));
 sky130_fd_sc_hd__a21oi_1 _09470_ (.A1(_03191_),
    .A2(_03755_),
    .B1(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__o21ai_0 _09471_ (.A1(_03189_),
    .A2(_03770_),
    .B1(_03799_),
    .Y(_00824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_220 ();
 sky130_fd_sc_hd__nor2_1 _09473_ (.A(_03201_),
    .B(_03750_),
    .Y(_03801_));
 sky130_fd_sc_hd__a21oi_1 _09474_ (.A1(net1517),
    .A2(_03750_),
    .B1(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nor2_1 _09475_ (.A(CPU_reset_a3),
    .B(_03802_),
    .Y(_00825_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(_03210_),
    .B(_03755_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(net1182),
    .B(_03750_),
    .Y(_03804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_219 ();
 sky130_fd_sc_hd__a21oi_1 _09479_ (.A1(_03803_),
    .A2(_03804_),
    .B1(net110),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _09480_ (.A(_03219_),
    .B(_03755_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(net1256),
    .B(_03750_),
    .Y(_03807_));
 sky130_fd_sc_hd__a21oi_1 _09482_ (.A1(_03806_),
    .A2(_03807_),
    .B1(CPU_reset_a3),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_03227_),
    .B(_03755_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(net1359),
    .B(_03750_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21oi_1 _09485_ (.A1(_03808_),
    .A2(_03809_),
    .B1(net109),
    .Y(_00828_));
 sky130_fd_sc_hd__nand3_1 _09486_ (.A(net1387),
    .B(net96),
    .C(_03750_),
    .Y(_03810_));
 sky130_fd_sc_hd__o31ai_1 _09487_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03750_),
    .B1(_03810_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand3_1 _09488_ (.A(net1400),
    .B(net96),
    .C(_03750_),
    .Y(_03811_));
 sky130_fd_sc_hd__o21ai_0 _09489_ (.A1(_03251_),
    .A2(_03750_),
    .B1(_03811_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand3_1 _09490_ (.A(net1392),
    .B(net96),
    .C(_03750_),
    .Y(_03812_));
 sky130_fd_sc_hd__o31ai_1 _09491_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03750_),
    .B1(_03812_),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2b_1 _09492_ (.A_N(\CPU_rd_a5[3] ),
    .B(\CPU_rd_a5[2] ),
    .Y(_03813_));
 sky130_fd_sc_hd__or3_1 _09493_ (.A(_02564_),
    .B(\CPU_rd_a3[3] ),
    .C(_01035_),
    .X(_03814_));
 sky130_fd_sc_hd__o21a_4 _09494_ (.A1(_01036_),
    .A2(_03813_),
    .B1(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__nor2_8 _09495_ (.A(_03361_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_8 _09496_ (.A(_02581_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_216 ();
 sky130_fd_sc_hd__o21ai_4 _09500_ (.A1(_01036_),
    .A2(_03813_),
    .B1(_03814_),
    .Y(_03821_));
 sky130_fd_sc_hd__nand2_8 _09501_ (.A(_03368_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_215 ();
 sky130_fd_sc_hd__and3_1 _09503_ (.A(net1832),
    .B(net97),
    .C(_03822_),
    .X(_03824_));
 sky130_fd_sc_hd__a21oi_1 _09504_ (.A1(_02588_),
    .A2(_03816_),
    .B1(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__o21ai_0 _09505_ (.A1(_02560_),
    .A2(_03817_),
    .B1(_03825_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_1 _09506_ (.A(_02636_),
    .B(_03816_),
    .Y(_03826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_214 ();
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(net1347),
    .B(_03822_),
    .Y(_03828_));
 sky130_fd_sc_hd__a21oi_1 _09509_ (.A1(_03826_),
    .A2(_03828_),
    .B1(net108),
    .Y(_00833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_213 ();
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(net1176),
    .B(_03822_),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _09512_ (.A(_02683_),
    .B(_03816_),
    .Y(_03831_));
 sky130_fd_sc_hd__a21oi_1 _09513_ (.A1(_03830_),
    .A2(_03831_),
    .B1(net109),
    .Y(_00834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_210 ();
 sky130_fd_sc_hd__nand3_1 _09517_ (.A(net1435),
    .B(net96),
    .C(_03822_),
    .Y(_03835_));
 sky130_fd_sc_hd__o21ai_0 _09518_ (.A1(_02713_),
    .A2(_03822_),
    .B1(_03835_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _09519_ (.A(_02748_),
    .B(_03816_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(net1131),
    .B(_03822_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21oi_1 _09521_ (.A1(_03836_),
    .A2(_03837_),
    .B1(net109),
    .Y(_00836_));
 sky130_fd_sc_hd__nand3_1 _09522_ (.A(net1428),
    .B(net97),
    .C(_03822_),
    .Y(_03838_));
 sky130_fd_sc_hd__o21ai_0 _09523_ (.A1(_02766_),
    .A2(_03822_),
    .B1(_03838_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand3_1 _09524_ (.A(net1369),
    .B(net97),
    .C(_03822_),
    .Y(_03839_));
 sky130_fd_sc_hd__o21ai_0 _09525_ (.A1(_02784_),
    .A2(_03822_),
    .B1(_03839_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand3_1 _09526_ (.A(net1417),
    .B(net97),
    .C(_03822_),
    .Y(_03840_));
 sky130_fd_sc_hd__o21ai_0 _09527_ (.A1(_02809_),
    .A2(_03822_),
    .B1(_03840_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand3_1 _09528_ (.A(net1526),
    .B(net97),
    .C(_03822_),
    .Y(_03841_));
 sky130_fd_sc_hd__o221ai_1 _09529_ (.A1(_02834_),
    .A2(_03822_),
    .B1(_03817_),
    .B2(_02832_),
    .C1(_03841_),
    .Y(_00840_));
 sky130_fd_sc_hd__and3_1 _09530_ (.A(net1731),
    .B(_02586_),
    .C(_03822_),
    .X(_03842_));
 sky130_fd_sc_hd__a31o_1 _09531_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03816_),
    .B1(_03842_),
    .X(_00841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_209 ();
 sky130_fd_sc_hd__and3_1 _09533_ (.A(net1769),
    .B(net97),
    .C(_03822_),
    .X(_03844_));
 sky130_fd_sc_hd__a21oi_1 _09534_ (.A1(_02884_),
    .A2(_03816_),
    .B1(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__o21ai_0 _09535_ (.A1(_02882_),
    .A2(_03817_),
    .B1(_03845_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_02889_),
    .B(_03822_),
    .Y(_03846_));
 sky130_fd_sc_hd__a21oi_1 _09537_ (.A1(net1650),
    .A2(_03822_),
    .B1(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__nor2_1 _09538_ (.A(net110),
    .B(_03847_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand3_1 _09539_ (.A(net1626),
    .B(net96),
    .C(_03822_),
    .Y(_03848_));
 sky130_fd_sc_hd__o221ai_1 _09540_ (.A1(_02909_),
    .A2(_03822_),
    .B1(_03817_),
    .B2(_02908_),
    .C1(_03848_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand3_1 _09541_ (.A(net1500),
    .B(_02586_),
    .C(_03822_),
    .Y(_03849_));
 sky130_fd_sc_hd__o221ai_1 _09542_ (.A1(_02936_),
    .A2(_03822_),
    .B1(_03817_),
    .B2(_02934_),
    .C1(_03849_),
    .Y(_00845_));
 sky130_fd_sc_hd__and3_1 _09543_ (.A(net1757),
    .B(_02586_),
    .C(_03822_),
    .X(_03850_));
 sky130_fd_sc_hd__a21oi_1 _09544_ (.A1(_02961_),
    .A2(_03816_),
    .B1(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__o21ai_0 _09545_ (.A1(_02959_),
    .A2(_03817_),
    .B1(_03851_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand3_1 _09546_ (.A(net1551),
    .B(_02586_),
    .C(_03822_),
    .Y(_03852_));
 sky130_fd_sc_hd__o221ai_1 _09547_ (.A1(_02984_),
    .A2(_03822_),
    .B1(_03817_),
    .B2(_02983_),
    .C1(_03852_),
    .Y(_00847_));
 sky130_fd_sc_hd__nand2_1 _09548_ (.A(net1290),
    .B(_03822_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_1 _09549_ (.A(_03009_),
    .B(_03816_),
    .Y(_03854_));
 sky130_fd_sc_hd__a21oi_1 _09550_ (.A1(_03853_),
    .A2(_03854_),
    .B1(net109),
    .Y(_00848_));
 sky130_fd_sc_hd__nor2_1 _09551_ (.A(_01035_),
    .B(_03822_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _09552_ (.A(_03031_),
    .B(_03816_),
    .Y(_03856_));
 sky130_fd_sc_hd__o21ai_0 _09553_ (.A1(net1712),
    .A2(_03816_),
    .B1(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__a311oi_1 _09554_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03855_),
    .B1(_03857_),
    .C1(net108),
    .Y(_00849_));
 sky130_fd_sc_hd__nand2_1 _09555_ (.A(_03053_),
    .B(_03816_),
    .Y(_03858_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(net1212),
    .B(_03822_),
    .Y(_03859_));
 sky130_fd_sc_hd__a21oi_1 _09557_ (.A1(_03858_),
    .A2(_03859_),
    .B1(net109),
    .Y(_00850_));
 sky130_fd_sc_hd__nand3_1 _09558_ (.A(net1518),
    .B(net97),
    .C(_03822_),
    .Y(_03860_));
 sky130_fd_sc_hd__o221ai_1 _09559_ (.A1(_03076_),
    .A2(_03822_),
    .B1(_03817_),
    .B2(_03074_),
    .C1(_03860_),
    .Y(_00851_));
 sky130_fd_sc_hd__and3_1 _09560_ (.A(net1764),
    .B(_02586_),
    .C(_03822_),
    .X(_03861_));
 sky130_fd_sc_hd__a21oi_1 _09561_ (.A1(_03100_),
    .A2(_03816_),
    .B1(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__o21ai_0 _09562_ (.A1(_03098_),
    .A2(_03817_),
    .B1(_03862_),
    .Y(_00852_));
 sky130_fd_sc_hd__a2111oi_0 _09563_ (.A1(net98),
    .A2(_03117_),
    .B1(_03822_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03863_));
 sky130_fd_sc_hd__nor2_1 _09564_ (.A(net1686),
    .B(_03816_),
    .Y(_03864_));
 sky130_fd_sc_hd__a2111oi_0 _09565_ (.A1(_03104_),
    .A2(_03816_),
    .B1(_03863_),
    .C1(_03864_),
    .D1(net108),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _09566_ (.A(net1410),
    .B(_03822_),
    .Y(_03865_));
 sky130_fd_sc_hd__o211ai_1 _09567_ (.A1(_03144_),
    .A2(_03822_),
    .B1(_03865_),
    .C1(_02586_),
    .Y(_00854_));
 sky130_fd_sc_hd__and3_1 _09568_ (.A(net1801),
    .B(_02586_),
    .C(_03822_),
    .X(_03866_));
 sky130_fd_sc_hd__a21oi_1 _09569_ (.A1(_03163_),
    .A2(_03816_),
    .B1(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__o21ai_0 _09570_ (.A1(_03161_),
    .A2(_03817_),
    .B1(_03867_),
    .Y(_00855_));
 sky130_fd_sc_hd__and3_1 _09571_ (.A(net1777),
    .B(net97),
    .C(_03822_),
    .X(_03868_));
 sky130_fd_sc_hd__a21oi_1 _09572_ (.A1(_03191_),
    .A2(_03816_),
    .B1(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o21ai_0 _09573_ (.A1(_03189_),
    .A2(_03817_),
    .B1(_03869_),
    .Y(_00856_));
 sky130_fd_sc_hd__nor2_1 _09574_ (.A(_03201_),
    .B(_03822_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_1 _09575_ (.A1(net1572),
    .A2(_03822_),
    .B1(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(CPU_reset_a3),
    .B(_03871_),
    .Y(_00857_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(_03210_),
    .B(_03816_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(net1168),
    .B(_03822_),
    .Y(_03873_));
 sky130_fd_sc_hd__a21oi_1 _09579_ (.A1(_03872_),
    .A2(_03873_),
    .B1(net110),
    .Y(_00858_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(_03219_),
    .B(_03816_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(net1451),
    .B(_03822_),
    .Y(_03875_));
 sky130_fd_sc_hd__a21oi_1 _09582_ (.A1(_03874_),
    .A2(_03875_),
    .B1(CPU_reset_a3),
    .Y(_00859_));
 sky130_fd_sc_hd__nand2_1 _09583_ (.A(_03227_),
    .B(_03816_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(net1295),
    .B(_03822_),
    .Y(_03877_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_208 ();
 sky130_fd_sc_hd__a21oi_1 _09586_ (.A1(_03876_),
    .A2(_03877_),
    .B1(net109),
    .Y(_00860_));
 sky130_fd_sc_hd__nand3_1 _09587_ (.A(net1423),
    .B(net96),
    .C(_03822_),
    .Y(_03879_));
 sky130_fd_sc_hd__o31ai_1 _09588_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03822_),
    .B1(_03879_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand3_1 _09589_ (.A(net1386),
    .B(net96),
    .C(_03822_),
    .Y(_03880_));
 sky130_fd_sc_hd__o21ai_0 _09590_ (.A1(_03251_),
    .A2(_03822_),
    .B1(_03880_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand3_1 _09591_ (.A(net1383),
    .B(net96),
    .C(_03822_),
    .Y(_03881_));
 sky130_fd_sc_hd__o31ai_1 _09592_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03822_),
    .B1(_03881_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand2_8 _09593_ (.A(_03431_),
    .B(_03821_),
    .Y(_03882_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_205 ();
 sky130_fd_sc_hd__a21oi_1 _09597_ (.A1(net1408),
    .A2(_03882_),
    .B1(CPU_reset_a3),
    .Y(_03886_));
 sky130_fd_sc_hd__o21ai_0 _09598_ (.A1(_03265_),
    .A2(_03882_),
    .B1(_03886_),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_8 _09599_ (.A(_03438_),
    .B(_03815_),
    .Y(_03887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_204 ();
 sky130_fd_sc_hd__nand2_1 _09601_ (.A(_02636_),
    .B(_03887_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(net1299),
    .B(_03882_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21oi_1 _09603_ (.A1(_03889_),
    .A2(_03890_),
    .B1(net108),
    .Y(_00865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_203 ();
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(net1284),
    .B(_03882_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(_02683_),
    .B(_03887_),
    .Y(_03893_));
 sky130_fd_sc_hd__a21oi_1 _09607_ (.A1(_03892_),
    .A2(_03893_),
    .B1(net109),
    .Y(_00866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_202 ();
 sky130_fd_sc_hd__nand3_1 _09609_ (.A(net1523),
    .B(net96),
    .C(_03882_),
    .Y(_03895_));
 sky130_fd_sc_hd__o21ai_0 _09610_ (.A1(_02713_),
    .A2(_03882_),
    .B1(_03895_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _09611_ (.A(_02748_),
    .B(_03887_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand2_1 _09612_ (.A(net1357),
    .B(_03882_),
    .Y(_03897_));
 sky130_fd_sc_hd__a21oi_1 _09613_ (.A1(_03896_),
    .A2(_03897_),
    .B1(net109),
    .Y(_00868_));
 sky130_fd_sc_hd__nand3_1 _09614_ (.A(net1373),
    .B(net97),
    .C(_03882_),
    .Y(_03898_));
 sky130_fd_sc_hd__o21ai_0 _09615_ (.A1(_02766_),
    .A2(_03882_),
    .B1(_03898_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand3_1 _09616_ (.A(net1643),
    .B(net97),
    .C(_03882_),
    .Y(_03899_));
 sky130_fd_sc_hd__o21ai_0 _09617_ (.A1(_02784_),
    .A2(_03882_),
    .B1(_03899_),
    .Y(_00870_));
 sky130_fd_sc_hd__nand3_1 _09618_ (.A(net1424),
    .B(net97),
    .C(_03882_),
    .Y(_03900_));
 sky130_fd_sc_hd__o21ai_0 _09619_ (.A1(_02809_),
    .A2(_03882_),
    .B1(_03900_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_8 _09620_ (.A(_02581_),
    .B(_03887_),
    .Y(_03901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_201 ();
 sky130_fd_sc_hd__nand3_1 _09622_ (.A(net1605),
    .B(net97),
    .C(_03882_),
    .Y(_03903_));
 sky130_fd_sc_hd__o221ai_1 _09623_ (.A1(_02834_),
    .A2(_03882_),
    .B1(_03901_),
    .B2(_02832_),
    .C1(_03903_),
    .Y(_00872_));
 sky130_fd_sc_hd__and3_1 _09624_ (.A(net1772),
    .B(_02586_),
    .C(_03882_),
    .X(_03904_));
 sky130_fd_sc_hd__a31o_1 _09625_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03887_),
    .B1(_03904_),
    .X(_00873_));
 sky130_fd_sc_hd__and3_1 _09626_ (.A(net1738),
    .B(net97),
    .C(_03882_),
    .X(_03905_));
 sky130_fd_sc_hd__a21oi_1 _09627_ (.A1(_02884_),
    .A2(_03887_),
    .B1(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__o21ai_0 _09628_ (.A1(_02882_),
    .A2(_03901_),
    .B1(_03906_),
    .Y(_00874_));
 sky130_fd_sc_hd__nor2_1 _09629_ (.A(_02889_),
    .B(_03882_),
    .Y(_03907_));
 sky130_fd_sc_hd__a21oi_1 _09630_ (.A1(net1659),
    .A2(_03882_),
    .B1(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__nor2_1 _09631_ (.A(CPU_reset_a3),
    .B(_03908_),
    .Y(_00875_));
 sky130_fd_sc_hd__nand3_1 _09632_ (.A(net1524),
    .B(net96),
    .C(_03882_),
    .Y(_03909_));
 sky130_fd_sc_hd__o221ai_1 _09633_ (.A1(_02909_),
    .A2(_03882_),
    .B1(_03901_),
    .B2(_02908_),
    .C1(_03909_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand3_1 _09634_ (.A(net1545),
    .B(_02586_),
    .C(_03882_),
    .Y(_03910_));
 sky130_fd_sc_hd__o221ai_1 _09635_ (.A1(_02936_),
    .A2(_03882_),
    .B1(_03901_),
    .B2(_02934_),
    .C1(_03910_),
    .Y(_00877_));
 sky130_fd_sc_hd__and3_1 _09636_ (.A(net1771),
    .B(_02586_),
    .C(_03882_),
    .X(_03911_));
 sky130_fd_sc_hd__a21oi_1 _09637_ (.A1(_02961_),
    .A2(_03887_),
    .B1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__o21ai_0 _09638_ (.A1(_02959_),
    .A2(_03901_),
    .B1(_03912_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand3_1 _09639_ (.A(net1617),
    .B(_02586_),
    .C(_03882_),
    .Y(_03913_));
 sky130_fd_sc_hd__o221ai_1 _09640_ (.A1(_02984_),
    .A2(_03882_),
    .B1(_03901_),
    .B2(_02983_),
    .C1(_03913_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_03009_),
    .B(_03887_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand2_1 _09642_ (.A(net1324),
    .B(_03882_),
    .Y(_03915_));
 sky130_fd_sc_hd__a21oi_1 _09643_ (.A1(_03914_),
    .A2(_03915_),
    .B1(net109),
    .Y(_00880_));
 sky130_fd_sc_hd__nor2_1 _09644_ (.A(_01035_),
    .B(_03882_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _09645_ (.A(_03031_),
    .B(_03887_),
    .Y(_03917_));
 sky130_fd_sc_hd__o21ai_0 _09646_ (.A1(net1705),
    .A2(_03887_),
    .B1(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a311oi_1 _09647_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03916_),
    .B1(_03918_),
    .C1(net108),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _09648_ (.A(_03053_),
    .B(_03887_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _09649_ (.A(net1354),
    .B(_03882_),
    .Y(_03920_));
 sky130_fd_sc_hd__a21oi_1 _09650_ (.A1(_03919_),
    .A2(_03920_),
    .B1(net109),
    .Y(_00882_));
 sky130_fd_sc_hd__nand3_1 _09651_ (.A(net1658),
    .B(_02586_),
    .C(_03882_),
    .Y(_03921_));
 sky130_fd_sc_hd__o221ai_1 _09652_ (.A1(_03076_),
    .A2(_03882_),
    .B1(_03901_),
    .B2(_03074_),
    .C1(_03921_),
    .Y(_00883_));
 sky130_fd_sc_hd__and3_1 _09653_ (.A(net1768),
    .B(net97),
    .C(_03882_),
    .X(_03922_));
 sky130_fd_sc_hd__a21oi_1 _09654_ (.A1(_03100_),
    .A2(_03887_),
    .B1(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__o21ai_0 _09655_ (.A1(_03098_),
    .A2(_03901_),
    .B1(_03923_),
    .Y(_00884_));
 sky130_fd_sc_hd__a2111oi_0 _09656_ (.A1(net98),
    .A2(_03117_),
    .B1(_03882_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03924_));
 sky130_fd_sc_hd__nor2_1 _09657_ (.A(net1619),
    .B(_03887_),
    .Y(_03925_));
 sky130_fd_sc_hd__a2111oi_0 _09658_ (.A1(_03104_),
    .A2(_03887_),
    .B1(_03924_),
    .C1(_03925_),
    .D1(net108),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _09659_ (.A(net1450),
    .B(_03882_),
    .Y(_03926_));
 sky130_fd_sc_hd__o211ai_1 _09660_ (.A1(_03144_),
    .A2(_03882_),
    .B1(_03926_),
    .C1(_02586_),
    .Y(_00886_));
 sky130_fd_sc_hd__and3_1 _09661_ (.A(net1810),
    .B(_02586_),
    .C(_03882_),
    .X(_03927_));
 sky130_fd_sc_hd__a21oi_1 _09662_ (.A1(_03163_),
    .A2(_03887_),
    .B1(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__o21ai_0 _09663_ (.A1(_03161_),
    .A2(_03901_),
    .B1(_03928_),
    .Y(_00887_));
 sky130_fd_sc_hd__and3_1 _09664_ (.A(net1734),
    .B(net97),
    .C(_03882_),
    .X(_03929_));
 sky130_fd_sc_hd__a21oi_1 _09665_ (.A1(_03191_),
    .A2(_03887_),
    .B1(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__o21ai_0 _09666_ (.A1(_03189_),
    .A2(_03901_),
    .B1(_03930_),
    .Y(_00888_));
 sky130_fd_sc_hd__nor2_1 _09667_ (.A(_03201_),
    .B(_03882_),
    .Y(_03931_));
 sky130_fd_sc_hd__a21oi_1 _09668_ (.A1(net1646),
    .A2(_03882_),
    .B1(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__nor2_1 _09669_ (.A(CPU_reset_a3),
    .B(_03932_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(_03210_),
    .B(_03887_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand2_1 _09671_ (.A(net1239),
    .B(_03882_),
    .Y(_03934_));
 sky130_fd_sc_hd__a21oi_1 _09672_ (.A1(_03933_),
    .A2(_03934_),
    .B1(net110),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _09673_ (.A(_03219_),
    .B(_03887_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(net1293),
    .B(_03882_),
    .Y(_03936_));
 sky130_fd_sc_hd__a21oi_1 _09675_ (.A1(_03935_),
    .A2(_03936_),
    .B1(CPU_reset_a3),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(_03227_),
    .B(_03887_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(net1233),
    .B(_03882_),
    .Y(_03938_));
 sky130_fd_sc_hd__a21oi_1 _09678_ (.A1(_03937_),
    .A2(_03938_),
    .B1(net109),
    .Y(_00892_));
 sky130_fd_sc_hd__nand3_1 _09679_ (.A(net1446),
    .B(net96),
    .C(_03882_),
    .Y(_03939_));
 sky130_fd_sc_hd__o31ai_1 _09680_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03882_),
    .B1(_03939_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand3_1 _09681_ (.A(net1448),
    .B(net96),
    .C(_03882_),
    .Y(_03940_));
 sky130_fd_sc_hd__o21ai_0 _09682_ (.A1(_03251_),
    .A2(_03882_),
    .B1(_03940_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3_1 _09683_ (.A(net1456),
    .B(net96),
    .C(_03882_),
    .Y(_03941_));
 sky130_fd_sc_hd__o31ai_1 _09684_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03882_),
    .B1(_03941_),
    .Y(_00895_));
 sky130_fd_sc_hd__nor2_8 _09685_ (.A(_02579_),
    .B(_03815_),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_8 _09686_ (.A(_02581_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_197 ();
 sky130_fd_sc_hd__nand2_8 _09691_ (.A(_02595_),
    .B(_03821_),
    .Y(_03948_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_196 ();
 sky130_fd_sc_hd__and3_1 _09693_ (.A(net1766),
    .B(net97),
    .C(_03948_),
    .X(_03950_));
 sky130_fd_sc_hd__a21oi_1 _09694_ (.A1(_02588_),
    .A2(_03942_),
    .B1(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__o21ai_0 _09695_ (.A1(_02560_),
    .A2(_03943_),
    .B1(_03951_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand2_1 _09696_ (.A(_02636_),
    .B(_03942_),
    .Y(_03952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_195 ();
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(net1385),
    .B(_03948_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21oi_1 _09699_ (.A1(_03952_),
    .A2(_03954_),
    .B1(net108),
    .Y(_00897_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_194 ();
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(net1389),
    .B(_03948_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand2_1 _09702_ (.A(_02683_),
    .B(_03942_),
    .Y(_03957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_193 ();
 sky130_fd_sc_hd__a21oi_1 _09704_ (.A1(_03956_),
    .A2(_03957_),
    .B1(net109),
    .Y(_00898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_190 ();
 sky130_fd_sc_hd__nand3_1 _09708_ (.A(net1487),
    .B(net96),
    .C(_03948_),
    .Y(_03962_));
 sky130_fd_sc_hd__o21ai_0 _09709_ (.A1(_02713_),
    .A2(_03948_),
    .B1(_03962_),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(_02748_),
    .B(_03942_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _09711_ (.A(net1457),
    .B(_03948_),
    .Y(_03964_));
 sky130_fd_sc_hd__a21oi_1 _09712_ (.A1(_03963_),
    .A2(_03964_),
    .B1(net109),
    .Y(_00900_));
 sky130_fd_sc_hd__nand3_1 _09713_ (.A(net1458),
    .B(net97),
    .C(_03948_),
    .Y(_03965_));
 sky130_fd_sc_hd__o21ai_0 _09714_ (.A1(_02766_),
    .A2(_03948_),
    .B1(_03965_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand3_1 _09715_ (.A(net1351),
    .B(net97),
    .C(_03948_),
    .Y(_03966_));
 sky130_fd_sc_hd__o21ai_0 _09716_ (.A1(_02784_),
    .A2(_03948_),
    .B1(_03966_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand3_1 _09717_ (.A(net1377),
    .B(net97),
    .C(_03948_),
    .Y(_03967_));
 sky130_fd_sc_hd__o21ai_0 _09718_ (.A1(_02809_),
    .A2(_03948_),
    .B1(_03967_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand3_1 _09719_ (.A(net1660),
    .B(net97),
    .C(_03948_),
    .Y(_03968_));
 sky130_fd_sc_hd__o221ai_1 _09720_ (.A1(_02834_),
    .A2(_03948_),
    .B1(_03943_),
    .B2(_02832_),
    .C1(_03968_),
    .Y(_00904_));
 sky130_fd_sc_hd__and3_1 _09721_ (.A(net1842),
    .B(_02586_),
    .C(_03948_),
    .X(_03969_));
 sky130_fd_sc_hd__a31o_1 _09722_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_03942_),
    .B1(_03969_),
    .X(_00905_));
 sky130_fd_sc_hd__and3_1 _09723_ (.A(net1746),
    .B(_02586_),
    .C(_03948_),
    .X(_03970_));
 sky130_fd_sc_hd__a21oi_1 _09724_ (.A1(_02884_),
    .A2(_03942_),
    .B1(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__o21ai_0 _09725_ (.A1(_02882_),
    .A2(_03943_),
    .B1(_03971_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(net1590),
    .B(_03948_),
    .Y(_03972_));
 sky130_fd_sc_hd__o211ai_1 _09727_ (.A1(_02889_),
    .A2(_03948_),
    .B1(_03972_),
    .C1(_02586_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand3_1 _09728_ (.A(net1554),
    .B(net96),
    .C(_03948_),
    .Y(_03973_));
 sky130_fd_sc_hd__o221ai_1 _09729_ (.A1(_02909_),
    .A2(_03948_),
    .B1(_03943_),
    .B2(_02908_),
    .C1(_03973_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand3_1 _09730_ (.A(net1672),
    .B(_02586_),
    .C(_03948_),
    .Y(_03974_));
 sky130_fd_sc_hd__o221ai_1 _09731_ (.A1(_02936_),
    .A2(_03948_),
    .B1(_03943_),
    .B2(_02934_),
    .C1(_03974_),
    .Y(_00909_));
 sky130_fd_sc_hd__and3_1 _09732_ (.A(net1841),
    .B(_02586_),
    .C(_03948_),
    .X(_03975_));
 sky130_fd_sc_hd__a21oi_1 _09733_ (.A1(_02961_),
    .A2(_03942_),
    .B1(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_0 _09734_ (.A1(_02959_),
    .A2(_03943_),
    .B1(_03976_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _09735_ (.A(net1516),
    .B(_02586_),
    .C(_03948_),
    .Y(_03977_));
 sky130_fd_sc_hd__o221ai_1 _09736_ (.A1(_02984_),
    .A2(_03948_),
    .B1(_03943_),
    .B2(_02983_),
    .C1(_03977_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _09737_ (.A(_03009_),
    .B(_03942_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(net1407),
    .B(_03948_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21oi_1 _09739_ (.A1(_03978_),
    .A2(_03979_),
    .B1(net109),
    .Y(_00912_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(_01035_),
    .B(_03948_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_03031_),
    .B(_03942_),
    .Y(_03981_));
 sky130_fd_sc_hd__o21ai_0 _09742_ (.A1(net1792),
    .A2(_03942_),
    .B1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__a311oi_1 _09743_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_03980_),
    .B1(_03982_),
    .C1(net108),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _09744_ (.A(_03053_),
    .B(_03942_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(net1433),
    .B(_03948_),
    .Y(_03984_));
 sky130_fd_sc_hd__a21oi_1 _09746_ (.A1(_03983_),
    .A2(_03984_),
    .B1(net109),
    .Y(_00914_));
 sky130_fd_sc_hd__nand3_1 _09747_ (.A(net1604),
    .B(net97),
    .C(_03948_),
    .Y(_03985_));
 sky130_fd_sc_hd__o221ai_1 _09748_ (.A1(_03076_),
    .A2(_03948_),
    .B1(_03943_),
    .B2(_03074_),
    .C1(_03985_),
    .Y(_00915_));
 sky130_fd_sc_hd__and3_1 _09749_ (.A(net1781),
    .B(_02586_),
    .C(_03948_),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_1 _09750_ (.A1(_03100_),
    .A2(_03942_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__o21ai_0 _09751_ (.A1(_03098_),
    .A2(_03943_),
    .B1(_03987_),
    .Y(_00916_));
 sky130_fd_sc_hd__a2111oi_0 _09752_ (.A1(net98),
    .A2(_03117_),
    .B1(_03948_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_03988_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(net1588),
    .B(_03942_),
    .Y(_03989_));
 sky130_fd_sc_hd__a2111oi_0 _09754_ (.A1(_03104_),
    .A2(_03942_),
    .B1(_03988_),
    .C1(_03989_),
    .D1(net108),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _09755_ (.A(net1449),
    .B(_03948_),
    .Y(_03990_));
 sky130_fd_sc_hd__o211ai_1 _09756_ (.A1(_03144_),
    .A2(_03948_),
    .B1(_03990_),
    .C1(net96),
    .Y(_00918_));
 sky130_fd_sc_hd__and3_1 _09757_ (.A(net1790),
    .B(_02586_),
    .C(_03948_),
    .X(_03991_));
 sky130_fd_sc_hd__a21oi_1 _09758_ (.A1(_03163_),
    .A2(_03942_),
    .B1(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__o21ai_0 _09759_ (.A1(_03161_),
    .A2(_03943_),
    .B1(_03992_),
    .Y(_00919_));
 sky130_fd_sc_hd__and3_1 _09760_ (.A(net1802),
    .B(net97),
    .C(_03948_),
    .X(_03993_));
 sky130_fd_sc_hd__a21oi_1 _09761_ (.A1(_03191_),
    .A2(_03942_),
    .B1(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__o21ai_0 _09762_ (.A1(_03189_),
    .A2(_03943_),
    .B1(_03994_),
    .Y(_00920_));
 sky130_fd_sc_hd__nor2_1 _09763_ (.A(_03201_),
    .B(_03948_),
    .Y(_03995_));
 sky130_fd_sc_hd__a21oi_1 _09764_ (.A1(net1668),
    .A2(_03948_),
    .B1(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__nor2_1 _09765_ (.A(CPU_reset_a3),
    .B(_03996_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_03210_),
    .B(_03942_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _09767_ (.A(net1243),
    .B(_03948_),
    .Y(_03998_));
 sky130_fd_sc_hd__a21oi_1 _09768_ (.A1(_03997_),
    .A2(_03998_),
    .B1(net110),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_03219_),
    .B(_03942_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(net1318),
    .B(_03948_),
    .Y(_04000_));
 sky130_fd_sc_hd__a21oi_1 _09771_ (.A1(_03999_),
    .A2(_04000_),
    .B1(CPU_reset_a3),
    .Y(_00923_));
 sky130_fd_sc_hd__nand2_1 _09772_ (.A(_03227_),
    .B(_03942_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(net1213),
    .B(_03948_),
    .Y(_04002_));
 sky130_fd_sc_hd__a21oi_1 _09774_ (.A1(_04001_),
    .A2(_04002_),
    .B1(net109),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _09775_ (.A(net1478),
    .B(net96),
    .C(_03948_),
    .Y(_04003_));
 sky130_fd_sc_hd__o31ai_1 _09776_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_03948_),
    .B1(_04003_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand3_1 _09777_ (.A(net1364),
    .B(net96),
    .C(_03948_),
    .Y(_04004_));
 sky130_fd_sc_hd__o21ai_0 _09778_ (.A1(_03251_),
    .A2(_03948_),
    .B1(_04004_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand3_1 _09779_ (.A(net1429),
    .B(net96),
    .C(_03948_),
    .Y(_04005_));
 sky130_fd_sc_hd__o31ai_1 _09780_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_03948_),
    .B1(_04005_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_8 _09781_ (.A(_03269_),
    .B(_03821_),
    .Y(_04006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_187 ();
 sky130_fd_sc_hd__nand2_1 _09785_ (.A(net1463),
    .B(_04006_),
    .Y(_04010_));
 sky130_fd_sc_hd__o211ai_1 _09786_ (.A1(_03265_),
    .A2(_04006_),
    .B1(_04010_),
    .C1(net96),
    .Y(_00928_));
 sky130_fd_sc_hd__nor2_8 _09787_ (.A(_03277_),
    .B(_03815_),
    .Y(_04011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_186 ();
 sky130_fd_sc_hd__nand2_1 _09789_ (.A(_02636_),
    .B(_04011_),
    .Y(_04013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_185 ();
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(net1253),
    .B(_04006_),
    .Y(_04015_));
 sky130_fd_sc_hd__a21oi_1 _09792_ (.A1(_04013_),
    .A2(_04015_),
    .B1(net108),
    .Y(_00929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_184 ();
 sky130_fd_sc_hd__nand2_1 _09794_ (.A(net1189),
    .B(_04006_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand2_1 _09795_ (.A(_02683_),
    .B(_04011_),
    .Y(_04018_));
 sky130_fd_sc_hd__a21oi_1 _09796_ (.A1(_04017_),
    .A2(_04018_),
    .B1(net109),
    .Y(_00930_));
 sky130_fd_sc_hd__nand3_1 _09797_ (.A(net1713),
    .B(net96),
    .C(_04006_),
    .Y(_04019_));
 sky130_fd_sc_hd__o21ai_0 _09798_ (.A1(_02713_),
    .A2(_04006_),
    .B1(_04019_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_02748_),
    .B(_04011_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_1 _09800_ (.A(net1298),
    .B(_04006_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21oi_1 _09801_ (.A1(_04020_),
    .A2(_04021_),
    .B1(net109),
    .Y(_00932_));
 sky130_fd_sc_hd__nand3_1 _09802_ (.A(net1445),
    .B(net97),
    .C(_04006_),
    .Y(_04022_));
 sky130_fd_sc_hd__o21ai_0 _09803_ (.A1(_02766_),
    .A2(_04006_),
    .B1(_04022_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand3_1 _09804_ (.A(net1379),
    .B(net97),
    .C(_04006_),
    .Y(_04023_));
 sky130_fd_sc_hd__o21ai_0 _09805_ (.A1(_02784_),
    .A2(_04006_),
    .B1(_04023_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _09806_ (.A(net1502),
    .B(net97),
    .C(_04006_),
    .Y(_04024_));
 sky130_fd_sc_hd__o21ai_0 _09807_ (.A1(_02809_),
    .A2(_04006_),
    .B1(_04024_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_8 _09808_ (.A(_02581_),
    .B(_04011_),
    .Y(_04025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_183 ();
 sky130_fd_sc_hd__nand3_1 _09810_ (.A(net1577),
    .B(net97),
    .C(_04006_),
    .Y(_04027_));
 sky130_fd_sc_hd__o221ai_1 _09811_ (.A1(_02834_),
    .A2(_04006_),
    .B1(_04025_),
    .B2(_02832_),
    .C1(_04027_),
    .Y(_00936_));
 sky130_fd_sc_hd__and3_1 _09812_ (.A(net1736),
    .B(_02586_),
    .C(_04006_),
    .X(_04028_));
 sky130_fd_sc_hd__a31o_1 _09813_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_04011_),
    .B1(_04028_),
    .X(_00937_));
 sky130_fd_sc_hd__and3_1 _09814_ (.A(net1750),
    .B(net97),
    .C(_04006_),
    .X(_04029_));
 sky130_fd_sc_hd__a21oi_1 _09815_ (.A1(_02884_),
    .A2(_04011_),
    .B1(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_0 _09816_ (.A1(_02882_),
    .A2(_04025_),
    .B1(_04030_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _09817_ (.A(net1537),
    .B(_04006_),
    .Y(_04031_));
 sky130_fd_sc_hd__o211ai_1 _09818_ (.A1(_02889_),
    .A2(_04006_),
    .B1(_04031_),
    .C1(net96),
    .Y(_00939_));
 sky130_fd_sc_hd__nand3_1 _09819_ (.A(net1540),
    .B(net96),
    .C(_04006_),
    .Y(_04032_));
 sky130_fd_sc_hd__o221ai_1 _09820_ (.A1(_02909_),
    .A2(_04006_),
    .B1(_04025_),
    .B2(_02908_),
    .C1(_04032_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand3_1 _09821_ (.A(net1489),
    .B(net96),
    .C(_04006_),
    .Y(_04033_));
 sky130_fd_sc_hd__o221ai_1 _09822_ (.A1(_02936_),
    .A2(_04006_),
    .B1(_04025_),
    .B2(_02934_),
    .C1(_04033_),
    .Y(_00941_));
 sky130_fd_sc_hd__and3_1 _09823_ (.A(net1828),
    .B(_02586_),
    .C(_04006_),
    .X(_04034_));
 sky130_fd_sc_hd__a21oi_1 _09824_ (.A1(_02961_),
    .A2(_04011_),
    .B1(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__o21ai_0 _09825_ (.A1(_02959_),
    .A2(_04025_),
    .B1(_04035_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand3_1 _09826_ (.A(net1510),
    .B(net97),
    .C(_04006_),
    .Y(_04036_));
 sky130_fd_sc_hd__o221ai_1 _09827_ (.A1(_02984_),
    .A2(_04006_),
    .B1(_04025_),
    .B2(_02983_),
    .C1(_04036_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _09828_ (.A(_03009_),
    .B(_04011_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(net1319),
    .B(_04006_),
    .Y(_04038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_182 ();
 sky130_fd_sc_hd__a21oi_1 _09831_ (.A1(_04037_),
    .A2(_04038_),
    .B1(net109),
    .Y(_00944_));
 sky130_fd_sc_hd__nor2_1 _09832_ (.A(_01035_),
    .B(_04006_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand2_1 _09833_ (.A(_03031_),
    .B(_04011_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_0 _09834_ (.A1(net1699),
    .A2(_04011_),
    .B1(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__a311oi_1 _09835_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_04040_),
    .B1(_04042_),
    .C1(net108),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(_03053_),
    .B(_04011_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(net1282),
    .B(_04006_),
    .Y(_04044_));
 sky130_fd_sc_hd__a21oi_1 _09838_ (.A1(_04043_),
    .A2(_04044_),
    .B1(net109),
    .Y(_00946_));
 sky130_fd_sc_hd__nand3_1 _09839_ (.A(net1565),
    .B(_02586_),
    .C(_04006_),
    .Y(_04045_));
 sky130_fd_sc_hd__o221ai_1 _09840_ (.A1(_03076_),
    .A2(_04006_),
    .B1(_04025_),
    .B2(_03074_),
    .C1(_04045_),
    .Y(_00947_));
 sky130_fd_sc_hd__and3_1 _09841_ (.A(net1812),
    .B(_02586_),
    .C(_04006_),
    .X(_04046_));
 sky130_fd_sc_hd__a21oi_1 _09842_ (.A1(_03100_),
    .A2(_04011_),
    .B1(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__o21ai_0 _09843_ (.A1(_03098_),
    .A2(_04025_),
    .B1(_04047_),
    .Y(_00948_));
 sky130_fd_sc_hd__a2111oi_0 _09844_ (.A1(net98),
    .A2(_03117_),
    .B1(_04006_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_04048_));
 sky130_fd_sc_hd__nor2_1 _09845_ (.A(net1508),
    .B(_04011_),
    .Y(_04049_));
 sky130_fd_sc_hd__a2111oi_0 _09846_ (.A1(_03104_),
    .A2(_04011_),
    .B1(_04048_),
    .C1(_04049_),
    .D1(net108),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(net1459),
    .B(_04006_),
    .Y(_04050_));
 sky130_fd_sc_hd__o211ai_1 _09848_ (.A1(_03144_),
    .A2(_04006_),
    .B1(_04050_),
    .C1(net96),
    .Y(_00950_));
 sky130_fd_sc_hd__and3_1 _09849_ (.A(net1793),
    .B(_02586_),
    .C(_04006_),
    .X(_04051_));
 sky130_fd_sc_hd__a21oi_1 _09850_ (.A1(_03163_),
    .A2(_04011_),
    .B1(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__o21ai_0 _09851_ (.A1(_03161_),
    .A2(_04025_),
    .B1(_04052_),
    .Y(_00951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_181 ();
 sky130_fd_sc_hd__and3_1 _09853_ (.A(net1765),
    .B(net97),
    .C(_04006_),
    .X(_04054_));
 sky130_fd_sc_hd__a21oi_1 _09854_ (.A1(_03191_),
    .A2(_04011_),
    .B1(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__o21ai_0 _09855_ (.A1(_03189_),
    .A2(_04025_),
    .B1(_04055_),
    .Y(_00952_));
 sky130_fd_sc_hd__nor2_1 _09856_ (.A(_03201_),
    .B(_04006_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21oi_1 _09857_ (.A1(net1530),
    .A2(_04006_),
    .B1(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nor2_1 _09858_ (.A(CPU_reset_a3),
    .B(_04057_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _09859_ (.A(_03210_),
    .B(_04011_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(net1338),
    .B(_04006_),
    .Y(_04059_));
 sky130_fd_sc_hd__a21oi_1 _09861_ (.A1(_04058_),
    .A2(_04059_),
    .B1(net110),
    .Y(_00954_));
 sky130_fd_sc_hd__nand2_1 _09862_ (.A(_03219_),
    .B(_04011_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(net1248),
    .B(_04006_),
    .Y(_04061_));
 sky130_fd_sc_hd__a21oi_1 _09864_ (.A1(_04060_),
    .A2(_04061_),
    .B1(CPU_reset_a3),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _09865_ (.A(_03227_),
    .B(_04011_),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(net1288),
    .B(_04006_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21oi_1 _09867_ (.A1(_04062_),
    .A2(_04063_),
    .B1(net110),
    .Y(_00956_));
 sky130_fd_sc_hd__nand3_1 _09868_ (.A(net1393),
    .B(net96),
    .C(_04006_),
    .Y(_04064_));
 sky130_fd_sc_hd__o31ai_1 _09869_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_04006_),
    .B1(_04064_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand3_1 _09870_ (.A(net1406),
    .B(net96),
    .C(_04006_),
    .Y(_04065_));
 sky130_fd_sc_hd__o21ai_0 _09871_ (.A1(_03251_),
    .A2(_04006_),
    .B1(_04065_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand3_1 _09872_ (.A(net1370),
    .B(net96),
    .C(_04006_),
    .Y(_04066_));
 sky130_fd_sc_hd__o31ai_1 _09873_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_04006_),
    .B1(_04066_),
    .Y(_00959_));
 sky130_fd_sc_hd__nor2_8 _09874_ (.A(_02567_),
    .B(_03361_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand2_8 _09875_ (.A(_02581_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_178 ();
 sky130_fd_sc_hd__nand2_8 _09879_ (.A(_02592_),
    .B(_03368_),
    .Y(_04072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_177 ();
 sky130_fd_sc_hd__and3_1 _09881_ (.A(net1840),
    .B(net97),
    .C(_04072_),
    .X(_04074_));
 sky130_fd_sc_hd__a21oi_1 _09882_ (.A1(_02588_),
    .A2(_04067_),
    .B1(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__o21ai_0 _09883_ (.A1(_02560_),
    .A2(_04068_),
    .B1(_04075_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_02636_),
    .B(_04067_),
    .Y(_04076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_176 ();
 sky130_fd_sc_hd__nand2_1 _09886_ (.A(net1185),
    .B(_04072_),
    .Y(_04078_));
 sky130_fd_sc_hd__a21oi_1 _09887_ (.A1(_04076_),
    .A2(_04078_),
    .B1(net108),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_1 _09888_ (.A(net1268),
    .B(_04072_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _09889_ (.A(_02683_),
    .B(_04067_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21oi_1 _09890_ (.A1(_04079_),
    .A2(_04080_),
    .B1(net109),
    .Y(_00962_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_172 ();
 sky130_fd_sc_hd__nand3_1 _09895_ (.A(net1501),
    .B(net96),
    .C(_04072_),
    .Y(_04085_));
 sky130_fd_sc_hd__o21ai_0 _09896_ (.A1(_02713_),
    .A2(_04072_),
    .B1(_04085_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(_02748_),
    .B(_04067_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_1 _09898_ (.A(net1184),
    .B(_04072_),
    .Y(_04087_));
 sky130_fd_sc_hd__a21oi_1 _09899_ (.A1(_04086_),
    .A2(_04087_),
    .B1(net109),
    .Y(_00964_));
 sky130_fd_sc_hd__nand3_1 _09900_ (.A(net1378),
    .B(net97),
    .C(_04072_),
    .Y(_04088_));
 sky130_fd_sc_hd__o21ai_0 _09901_ (.A1(_02766_),
    .A2(_04072_),
    .B1(_04088_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand3_1 _09902_ (.A(net1470),
    .B(net97),
    .C(_04072_),
    .Y(_04089_));
 sky130_fd_sc_hd__o21ai_0 _09903_ (.A1(_02784_),
    .A2(_04072_),
    .B1(_04089_),
    .Y(_00966_));
 sky130_fd_sc_hd__nand3_1 _09904_ (.A(net1452),
    .B(net97),
    .C(_04072_),
    .Y(_04090_));
 sky130_fd_sc_hd__o21ai_0 _09905_ (.A1(_02809_),
    .A2(_04072_),
    .B1(_04090_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand3_1 _09906_ (.A(net1595),
    .B(net97),
    .C(_04072_),
    .Y(_04091_));
 sky130_fd_sc_hd__o221ai_1 _09907_ (.A1(_02834_),
    .A2(_04072_),
    .B1(_04068_),
    .B2(_02832_),
    .C1(_04091_),
    .Y(_00968_));
 sky130_fd_sc_hd__and3_1 _09908_ (.A(net1776),
    .B(_02586_),
    .C(_04072_),
    .X(_04092_));
 sky130_fd_sc_hd__a31o_1 _09909_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_04067_),
    .B1(_04092_),
    .X(_00969_));
 sky130_fd_sc_hd__and3_1 _09910_ (.A(net1735),
    .B(net97),
    .C(_04072_),
    .X(_04093_));
 sky130_fd_sc_hd__a21oi_1 _09911_ (.A1(_02884_),
    .A2(_04067_),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__o21ai_0 _09912_ (.A1(_02882_),
    .A2(_04068_),
    .B1(_04094_),
    .Y(_00970_));
 sky130_fd_sc_hd__nor2_1 _09913_ (.A(_02889_),
    .B(_04072_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_1 _09914_ (.A1(net1521),
    .A2(_04072_),
    .B1(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__nor2_1 _09915_ (.A(CPU_reset_a3),
    .B(_04096_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand3_1 _09916_ (.A(net1538),
    .B(net96),
    .C(_04072_),
    .Y(_04097_));
 sky130_fd_sc_hd__o221ai_1 _09917_ (.A1(_02909_),
    .A2(_04072_),
    .B1(_04068_),
    .B2(_02908_),
    .C1(_04097_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand3_1 _09918_ (.A(net1480),
    .B(_02586_),
    .C(_04072_),
    .Y(_04098_));
 sky130_fd_sc_hd__o221ai_1 _09919_ (.A1(_02936_),
    .A2(_04072_),
    .B1(_04068_),
    .B2(_02934_),
    .C1(_04098_),
    .Y(_00973_));
 sky130_fd_sc_hd__and3_1 _09920_ (.A(net1778),
    .B(_02586_),
    .C(_04072_),
    .X(_04099_));
 sky130_fd_sc_hd__a21oi_1 _09921_ (.A1(_02961_),
    .A2(_04067_),
    .B1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__o21ai_0 _09922_ (.A1(_02959_),
    .A2(_04068_),
    .B1(_04100_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_1 _09923_ (.A(net1584),
    .B(_02586_),
    .C(_04072_),
    .Y(_04101_));
 sky130_fd_sc_hd__o221ai_1 _09924_ (.A1(_02984_),
    .A2(_04072_),
    .B1(_04068_),
    .B2(_02983_),
    .C1(_04101_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _09925_ (.A(_03009_),
    .B(_04067_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_1 _09926_ (.A(net1331),
    .B(_04072_),
    .Y(_04103_));
 sky130_fd_sc_hd__a21oi_1 _09927_ (.A1(_04102_),
    .A2(_04103_),
    .B1(net109),
    .Y(_00976_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(_01035_),
    .B(_04072_),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _09929_ (.A(_03031_),
    .B(_04067_),
    .Y(_04105_));
 sky130_fd_sc_hd__o21ai_0 _09930_ (.A1(net1701),
    .A2(_04067_),
    .B1(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a311oi_1 _09931_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_04104_),
    .B1(_04106_),
    .C1(net108),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_1 _09932_ (.A(_03053_),
    .B(_04067_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(net1270),
    .B(_04072_),
    .Y(_04108_));
 sky130_fd_sc_hd__a21oi_1 _09934_ (.A1(_04107_),
    .A2(_04108_),
    .B1(net109),
    .Y(_00978_));
 sky130_fd_sc_hd__nand3_1 _09935_ (.A(net1495),
    .B(_02586_),
    .C(_04072_),
    .Y(_04109_));
 sky130_fd_sc_hd__o221ai_1 _09936_ (.A1(_03076_),
    .A2(_04072_),
    .B1(_04068_),
    .B2(_03074_),
    .C1(_04109_),
    .Y(_00979_));
 sky130_fd_sc_hd__and3_1 _09937_ (.A(net1733),
    .B(_02586_),
    .C(_04072_),
    .X(_04110_));
 sky130_fd_sc_hd__a21oi_1 _09938_ (.A1(_03100_),
    .A2(_04067_),
    .B1(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__o21ai_0 _09939_ (.A1(_03098_),
    .A2(_04068_),
    .B1(_04111_),
    .Y(_00980_));
 sky130_fd_sc_hd__a2111oi_0 _09940_ (.A1(net98),
    .A2(_03117_),
    .B1(_04072_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _09941_ (.A(net1547),
    .B(_04067_),
    .Y(_04113_));
 sky130_fd_sc_hd__a2111oi_0 _09942_ (.A1(_03104_),
    .A2(_04067_),
    .B1(_04112_),
    .C1(_04113_),
    .D1(net108),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _09943_ (.A(_03144_),
    .B(_04072_),
    .Y(_04114_));
 sky130_fd_sc_hd__a21oi_1 _09944_ (.A1(net1663),
    .A2(_04072_),
    .B1(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__nor2_1 _09945_ (.A(net110),
    .B(_04115_),
    .Y(_00982_));
 sky130_fd_sc_hd__and3_1 _09946_ (.A(net1774),
    .B(_02586_),
    .C(_04072_),
    .X(_04116_));
 sky130_fd_sc_hd__a21oi_1 _09947_ (.A1(_03163_),
    .A2(_04067_),
    .B1(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__o21ai_0 _09948_ (.A1(_03161_),
    .A2(_04068_),
    .B1(_04117_),
    .Y(_00983_));
 sky130_fd_sc_hd__and3_1 _09949_ (.A(net1780),
    .B(net97),
    .C(_04072_),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_1 _09950_ (.A1(_03191_),
    .A2(_04067_),
    .B1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__o21ai_0 _09951_ (.A1(_03189_),
    .A2(_04068_),
    .B1(_04119_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _09952_ (.A(net1486),
    .B(_04072_),
    .Y(_04120_));
 sky130_fd_sc_hd__o211ai_1 _09953_ (.A1(_03201_),
    .A2(_04072_),
    .B1(_04120_),
    .C1(net96),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _09954_ (.A(_03210_),
    .B(_04067_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(net1149),
    .B(_04072_),
    .Y(_04122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_171 ();
 sky130_fd_sc_hd__a21oi_1 _09957_ (.A1(_04121_),
    .A2(_04122_),
    .B1(net110),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _09958_ (.A(_03219_),
    .B(_04067_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _09959_ (.A(net1325),
    .B(_04072_),
    .Y(_04125_));
 sky130_fd_sc_hd__a21oi_1 _09960_ (.A1(_04124_),
    .A2(_04125_),
    .B1(CPU_reset_a3),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _09961_ (.A(_03227_),
    .B(_04067_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(net1343),
    .B(_04072_),
    .Y(_04127_));
 sky130_fd_sc_hd__a21oi_1 _09963_ (.A1(_04126_),
    .A2(_04127_),
    .B1(net109),
    .Y(_00988_));
 sky130_fd_sc_hd__nand3_1 _09964_ (.A(net1464),
    .B(net96),
    .C(_04072_),
    .Y(_04128_));
 sky130_fd_sc_hd__o31ai_1 _09965_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_04072_),
    .B1(_04128_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand3_1 _09966_ (.A(net1425),
    .B(net96),
    .C(_04072_),
    .Y(_04129_));
 sky130_fd_sc_hd__o21ai_0 _09967_ (.A1(_03251_),
    .A2(_04072_),
    .B1(_04129_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand3_1 _09968_ (.A(net1374),
    .B(net96),
    .C(_04072_),
    .Y(_04130_));
 sky130_fd_sc_hd__o31ai_1 _09969_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_04072_),
    .B1(_04130_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_8 _09970_ (.A(_02592_),
    .B(_03431_),
    .Y(_04131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_168 ();
 sky130_fd_sc_hd__a21oi_1 _09974_ (.A1(net1514),
    .A2(_04131_),
    .B1(net108),
    .Y(_04135_));
 sky130_fd_sc_hd__o21ai_0 _09975_ (.A1(_03265_),
    .A2(_04131_),
    .B1(_04135_),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_8 _09976_ (.A(_02567_),
    .B(_03438_),
    .Y(_04136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_167 ();
 sky130_fd_sc_hd__nand2_1 _09978_ (.A(_02636_),
    .B(_04136_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _09979_ (.A(net1366),
    .B(_04131_),
    .Y(_04139_));
 sky130_fd_sc_hd__a21oi_1 _09980_ (.A1(_04138_),
    .A2(_04139_),
    .B1(net108),
    .Y(_00993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_166 ();
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(net1358),
    .B(_04131_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _09983_ (.A(_02683_),
    .B(_04136_),
    .Y(_04142_));
 sky130_fd_sc_hd__a21oi_1 _09984_ (.A1(_04141_),
    .A2(_04142_),
    .B1(net109),
    .Y(_00994_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__nand3_1 _09986_ (.A(net1415),
    .B(net96),
    .C(_04131_),
    .Y(_04144_));
 sky130_fd_sc_hd__o21ai_0 _09987_ (.A1(_02713_),
    .A2(_04131_),
    .B1(_04144_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _09988_ (.A(_02748_),
    .B(_04136_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(net1177),
    .B(_04131_),
    .Y(_04146_));
 sky130_fd_sc_hd__a21oi_1 _09990_ (.A1(_04145_),
    .A2(_04146_),
    .B1(net109),
    .Y(_00996_));
 sky130_fd_sc_hd__nand3_1 _09991_ (.A(net1365),
    .B(net97),
    .C(_04131_),
    .Y(_04147_));
 sky130_fd_sc_hd__o21ai_0 _09992_ (.A1(_02766_),
    .A2(_04131_),
    .B1(_04147_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand3_1 _09993_ (.A(net1395),
    .B(net97),
    .C(_04131_),
    .Y(_04148_));
 sky130_fd_sc_hd__o21ai_0 _09994_ (.A1(_02784_),
    .A2(_04131_),
    .B1(_04148_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand3_1 _09995_ (.A(net1390),
    .B(net97),
    .C(_04131_),
    .Y(_04149_));
 sky130_fd_sc_hd__o21ai_0 _09996_ (.A1(_02809_),
    .A2(_04131_),
    .B1(_04149_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_8 _09997_ (.A(_02581_),
    .B(_04136_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand3_1 _09998_ (.A(net1543),
    .B(net97),
    .C(_04131_),
    .Y(_04151_));
 sky130_fd_sc_hd__o221ai_1 _09999_ (.A1(_02834_),
    .A2(_04131_),
    .B1(_04150_),
    .B2(_02832_),
    .C1(_04151_),
    .Y(_01000_));
 sky130_fd_sc_hd__and3_1 _10000_ (.A(net1836),
    .B(_02586_),
    .C(_04131_),
    .X(_04152_));
 sky130_fd_sc_hd__a31o_1 _10001_ (.A1(_02854_),
    .A2(_02856_),
    .A3(_04136_),
    .B1(_04152_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _10002_ (.A(net1791),
    .B(net97),
    .C(_04131_),
    .X(_04153_));
 sky130_fd_sc_hd__a21oi_1 _10003_ (.A1(_02884_),
    .A2(_04136_),
    .B1(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__o21ai_0 _10004_ (.A1(_02882_),
    .A2(_04150_),
    .B1(_04154_),
    .Y(_01002_));
 sky130_fd_sc_hd__nor2_1 _10005_ (.A(_02889_),
    .B(_04131_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21oi_1 _10006_ (.A1(net1609),
    .A2(_04131_),
    .B1(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nor2_1 _10007_ (.A(CPU_reset_a3),
    .B(_04156_),
    .Y(_01003_));
 sky130_fd_sc_hd__nand3_1 _10008_ (.A(net1656),
    .B(net97),
    .C(_04131_),
    .Y(_04157_));
 sky130_fd_sc_hd__o221ai_1 _10009_ (.A1(_02909_),
    .A2(_04131_),
    .B1(_04150_),
    .B2(_02908_),
    .C1(_04157_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand3_1 _10010_ (.A(net1616),
    .B(_02586_),
    .C(_04131_),
    .Y(_04158_));
 sky130_fd_sc_hd__o221ai_1 _10011_ (.A1(_02936_),
    .A2(_04131_),
    .B1(_04150_),
    .B2(_02934_),
    .C1(_04158_),
    .Y(_01005_));
 sky130_fd_sc_hd__and3_1 _10012_ (.A(net1740),
    .B(_02586_),
    .C(_04131_),
    .X(_04159_));
 sky130_fd_sc_hd__a21oi_1 _10013_ (.A1(_02961_),
    .A2(_04136_),
    .B1(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__o21ai_0 _10014_ (.A1(_02959_),
    .A2(_04150_),
    .B1(_04160_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand3_1 _10015_ (.A(net1600),
    .B(_02586_),
    .C(_04131_),
    .Y(_04161_));
 sky130_fd_sc_hd__o221ai_1 _10016_ (.A1(_02984_),
    .A2(_04131_),
    .B1(_04150_),
    .B2(_02983_),
    .C1(_04161_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _10017_ (.A(_03009_),
    .B(_04136_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(net1375),
    .B(_04131_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_1 _10019_ (.A1(_04162_),
    .A2(_04163_),
    .B1(net109),
    .Y(_01008_));
 sky130_fd_sc_hd__nor2_1 _10020_ (.A(_01035_),
    .B(_04131_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_03031_),
    .B(_04136_),
    .Y(_04165_));
 sky130_fd_sc_hd__o21ai_0 _10022_ (.A1(net1711),
    .A2(_04136_),
    .B1(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__a311oi_1 _10023_ (.A1(_03018_),
    .A2(_03026_),
    .A3(_04164_),
    .B1(_04166_),
    .C1(net108),
    .Y(_01009_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(net1346),
    .B(_04131_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand2_1 _10025_ (.A(_03053_),
    .B(_04136_),
    .Y(_04168_));
 sky130_fd_sc_hd__a21oi_1 _10026_ (.A1(_04167_),
    .A2(_04168_),
    .B1(net109),
    .Y(_01010_));
 sky130_fd_sc_hd__nand3_1 _10027_ (.A(net1651),
    .B(_02586_),
    .C(_04131_),
    .Y(_04169_));
 sky130_fd_sc_hd__o221ai_1 _10028_ (.A1(_03076_),
    .A2(_04131_),
    .B1(_04150_),
    .B2(_03074_),
    .C1(_04169_),
    .Y(_01011_));
 sky130_fd_sc_hd__and3_1 _10029_ (.A(net1726),
    .B(net97),
    .C(_04131_),
    .X(_04170_));
 sky130_fd_sc_hd__a21oi_1 _10030_ (.A1(_03100_),
    .A2(_04136_),
    .B1(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__o21ai_0 _10031_ (.A1(_03098_),
    .A2(_04150_),
    .B1(_04171_),
    .Y(_01012_));
 sky130_fd_sc_hd__a2111oi_0 _10032_ (.A1(net98),
    .A2(_03117_),
    .B1(_04131_),
    .C1(_03135_),
    .D1(_01035_),
    .Y(_04172_));
 sky130_fd_sc_hd__nor2_1 _10033_ (.A(net1528),
    .B(_04136_),
    .Y(_04173_));
 sky130_fd_sc_hd__a2111oi_0 _10034_ (.A1(_03104_),
    .A2(_04136_),
    .B1(_04172_),
    .C1(_04173_),
    .D1(net108),
    .Y(_01013_));
 sky130_fd_sc_hd__nor2_1 _10035_ (.A(_03144_),
    .B(_04131_),
    .Y(_04174_));
 sky130_fd_sc_hd__a21oi_1 _10036_ (.A1(net1570),
    .A2(_04131_),
    .B1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nor2_1 _10037_ (.A(net110),
    .B(_04175_),
    .Y(_01014_));
 sky130_fd_sc_hd__and3_1 _10038_ (.A(net1739),
    .B(_02586_),
    .C(_04131_),
    .X(_04176_));
 sky130_fd_sc_hd__a21oi_1 _10039_ (.A1(_03163_),
    .A2(_04136_),
    .B1(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__o21ai_0 _10040_ (.A1(_03161_),
    .A2(_04150_),
    .B1(_04177_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _10041_ (.A(net1805),
    .B(net97),
    .C(_04131_),
    .X(_04178_));
 sky130_fd_sc_hd__a21oi_1 _10042_ (.A1(_03191_),
    .A2(_04136_),
    .B1(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__o21ai_0 _10043_ (.A1(_03189_),
    .A2(_04150_),
    .B1(_04179_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(net1474),
    .B(_04131_),
    .Y(_04180_));
 sky130_fd_sc_hd__o211ai_1 _10045_ (.A1(_03201_),
    .A2(_04131_),
    .B1(_04180_),
    .C1(net96),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_03210_),
    .B(_04136_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _10047_ (.A(net1327),
    .B(_04131_),
    .Y(_04182_));
 sky130_fd_sc_hd__a21oi_1 _10048_ (.A1(_04181_),
    .A2(_04182_),
    .B1(net110),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _10049_ (.A(_03219_),
    .B(_04136_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _10050_ (.A(net1388),
    .B(_04131_),
    .Y(_04184_));
 sky130_fd_sc_hd__a21oi_1 _10051_ (.A1(_04183_),
    .A2(_04184_),
    .B1(CPU_reset_a3),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _10052_ (.A(_03227_),
    .B(_04136_),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(net1103),
    .B(_04131_),
    .Y(_04186_));
 sky130_fd_sc_hd__a21oi_1 _10054_ (.A1(_04185_),
    .A2(_04186_),
    .B1(net110),
    .Y(_01020_));
 sky130_fd_sc_hd__nand3_1 _10055_ (.A(net1430),
    .B(net96),
    .C(_04131_),
    .Y(_04187_));
 sky130_fd_sc_hd__o31ai_1 _10056_ (.A1(_03236_),
    .A2(_03238_),
    .A3(_04131_),
    .B1(_04187_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand3_1 _10057_ (.A(net1350),
    .B(net96),
    .C(_04131_),
    .Y(_04188_));
 sky130_fd_sc_hd__o21ai_0 _10058_ (.A1(_03251_),
    .A2(_04131_),
    .B1(_04188_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand3_1 _10059_ (.A(net1432),
    .B(net96),
    .C(_04131_),
    .Y(_04189_));
 sky130_fd_sc_hd__o31ai_1 _10060_ (.A1(_03259_),
    .A2(_03261_),
    .A3(_04131_),
    .B1(_04189_),
    .Y(_01023_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(\CPU_inc_pc_a3[2] ),
    .B(_01119_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21oi_1 _10062_ (.A1(net192),
    .A2(_01119_),
    .B1(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__mux2i_1 _10063_ (.A0(net1302),
    .A1(_04191_),
    .S(_01118_),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2_1 _10064_ (.A(net1214),
    .B(net1303),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _10065_ (.A(net1016),
    .B(CPU_valid_load_a3),
    .Y(_04193_));
 sky130_fd_sc_hd__nand2_1 _10066_ (.A(\CPU_inc_pc_a1[3] ),
    .B(_01119_),
    .Y(_04194_));
 sky130_fd_sc_hd__nor2_1 _10067_ (.A(\CPU_br_tgt_pc_a3[3] ),
    .B(_01118_),
    .Y(_04195_));
 sky130_fd_sc_hd__a311oi_1 _10068_ (.A1(_01118_),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04195_),
    .C1(CPU_reset_a1),
    .Y(_01025_));
 sky130_fd_sc_hd__mux2i_1 _10069_ (.A0(net1556),
    .A1(\CPU_inc_pc_a1[4] ),
    .S(_01119_),
    .Y(_04196_));
 sky130_fd_sc_hd__or3b_1 _10070_ (.A(net1214),
    .B(_01118_),
    .C_N(\CPU_br_tgt_pc_a3[4] ),
    .X(_04197_));
 sky130_fd_sc_hd__o31ai_1 _10071_ (.A1(net1214),
    .A2(CPU_valid_taken_br_a3),
    .A3(net1557),
    .B1(_04197_),
    .Y(_01026_));
 sky130_fd_sc_hd__mux2i_1 _10072_ (.A0(net1581),
    .A1(\CPU_inc_pc_a1[5] ),
    .S(_01119_),
    .Y(_04198_));
 sky130_fd_sc_hd__or3b_1 _10073_ (.A(net1214),
    .B(_01118_),
    .C_N(\CPU_br_tgt_pc_a3[5] ),
    .X(_04199_));
 sky130_fd_sc_hd__o31ai_1 _10074_ (.A1(net1214),
    .A2(CPU_valid_taken_br_a3),
    .A3(net1582),
    .B1(_04199_),
    .Y(_01027_));
 sky130_fd_sc_hd__nor4_1 _10075_ (.A(_05822_),
    .B(_05817_),
    .C(_05820_),
    .D(_01122_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _10076_ (.A(net751),
    .B(CPU_valid_load_a3),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(net138),
    .B(_01119_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_1 _10078_ (.A(\CPU_br_tgt_pc_a3[0] ),
    .B(_01118_),
    .Y(_04202_));
 sky130_fd_sc_hd__a311oi_1 _10079_ (.A1(_01118_),
    .A2(_04200_),
    .A3(_04201_),
    .B1(_04202_),
    .C1(CPU_reset_a1),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _10080_ (.A(net1030),
    .B(CPU_valid_load_a3),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _10081_ (.A(net148),
    .B(_01119_),
    .Y(_04204_));
 sky130_fd_sc_hd__nor2_1 _10082_ (.A(\CPU_br_tgt_pc_a3[1] ),
    .B(_01118_),
    .Y(_04205_));
 sky130_fd_sc_hd__a311oi_1 _10083_ (.A1(_01118_),
    .A2(_04203_),
    .A3(_04204_),
    .B1(_04205_),
    .C1(CPU_reset_a1),
    .Y(_01030_));
 sky130_fd_sc_hd__nor3_1 _10084_ (.A(_05818_),
    .B(_05817_),
    .C(_05820_),
    .Y(_04206_));
 sky130_fd_sc_hd__nor2_1 _10085_ (.A(_01147_),
    .B(_04206_),
    .Y(_01031_));
 sky130_fd_sc_hd__nor2_1 _10086_ (.A(net827),
    .B(_01138_),
    .Y(_04207_));
 sky130_fd_sc_hd__nor2_1 _10087_ (.A(_05822_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_1 _10088_ (.A(net1291),
    .B(_04208_),
    .Y(_01032_));
 sky130_fd_sc_hd__a21oi_1 _10089_ (.A1(_01130_),
    .A2(_01149_),
    .B1(_01147_),
    .Y(_01033_));
 sky130_fd_sc_hd__nor2_1 _10090_ (.A(net1291),
    .B(_01132_),
    .Y(_01034_));
 sky130_fd_sc_hd__xnor2_1 _10091_ (.A(_05522_),
    .B(_05810_),
    .Y(\CPU_br_tgt_pc_a2[2] ));
 sky130_fd_sc_hd__a21o_1 _10092_ (.A1(_05815_),
    .A2(_05808_),
    .B1(_05807_),
    .X(_04209_));
 sky130_fd_sc_hd__a21oi_1 _10093_ (.A1(_05810_),
    .A2(_04209_),
    .B1(_05809_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _10094_ (.A(_05812_),
    .B(_04210_),
    .Y(\CPU_br_tgt_pc_a2[3] ));
 sky130_fd_sc_hd__inv_1 _10095_ (.A(_05522_),
    .Y(_04211_));
 sky130_fd_sc_hd__a21o_1 _10096_ (.A1(_04211_),
    .A2(_05810_),
    .B1(_05809_),
    .X(_04212_));
 sky130_fd_sc_hd__a21oi_1 _10097_ (.A1(_05812_),
    .A2(_04212_),
    .B1(_05811_),
    .Y(_04213_));
 sky130_fd_sc_hd__xnor2_1 _10098_ (.A(_05814_),
    .B(_04213_),
    .Y(\CPU_br_tgt_pc_a2[4] ));
 sky130_fd_sc_hd__xor2_1 _10099_ (.A(net1693),
    .B(net179),
    .X(_04214_));
 sky130_fd_sc_hd__inv_1 _10100_ (.A(_05812_),
    .Y(_04215_));
 sky130_fd_sc_hd__o21bai_1 _10101_ (.A1(_04215_),
    .A2(_04210_),
    .B1_N(_05811_),
    .Y(_04216_));
 sky130_fd_sc_hd__a21oi_1 _10102_ (.A1(_05814_),
    .A2(_04216_),
    .B1(_05813_),
    .Y(_04217_));
 sky130_fd_sc_hd__xnor2_1 _10103_ (.A(_04214_),
    .B(_04217_),
    .Y(\CPU_br_tgt_pc_a2[5] ));
 sky130_fd_sc_hd__nor2_1 _10104_ (.A(_01129_),
    .B(_01147_),
    .Y(\CPU_imem_rd_data_a1[20] ));
 sky130_fd_sc_hd__nand2_1 _10105_ (.A(_01121_),
    .B(_01146_),
    .Y(_04218_));
 sky130_fd_sc_hd__o21ai_1 _10106_ (.A1(_01140_),
    .A2(_01153_),
    .B1(_04218_),
    .Y(\CPU_imm_a1[0] ));
 sky130_fd_sc_hd__nor4_1 _10107_ (.A(_05822_),
    .B(_05817_),
    .C(_05820_),
    .D(_01122_),
    .Y(\CPU_imm_a1[11] ));
 sky130_fd_sc_hd__mux2i_1 _10108_ (.A0(_05818_),
    .A1(_05817_),
    .S(\CPU_imem_rd_addr_a1[3] ),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_1 _10109_ (.A(_05817_),
    .B(_01121_),
    .Y(_04220_));
 sky130_fd_sc_hd__o21ai_0 _10110_ (.A1(net1569),
    .A2(_04219_),
    .B1(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__and2_0 _10111_ (.A(_01133_),
    .B(_04221_),
    .X(\CPU_imem_rd_data_a1[21] ));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(_01148_),
    .B(\CPU_imem_rd_data_a1[21] ),
    .Y(_04222_));
 sky130_fd_sc_hd__o21ai_0 _10113_ (.A1(_01140_),
    .A2(_01153_),
    .B1(_04222_),
    .Y(\CPU_imm_a1[1] ));
 sky130_fd_sc_hd__a31oi_1 _10114_ (.A1(_01120_),
    .A2(net1833),
    .A3(_05820_),
    .B1(\CPU_dec_bits_a1[10] ),
    .Y(_04223_));
 sky130_fd_sc_hd__a21boi_0 _10115_ (.A1(_04220_),
    .A2(_04223_),
    .B1_N(_01133_),
    .Y(\CPU_imem_rd_data_a1[22] ));
 sky130_fd_sc_hd__and2_0 _10116_ (.A(_01148_),
    .B(\CPU_imem_rd_data_a1[22] ),
    .X(CPU_is_load_a1));
 sky130_fd_sc_hd__or2_0 _10117_ (.A(CPU_is_s_instr_a1),
    .B(CPU_is_load_a1),
    .X(\CPU_imm_a1[2] ));
 sky130_fd_sc_hd__or2_0 _10118_ (.A(\CPU_dec_bits_a1[10] ),
    .B(\CPU_imem_rd_data_a1[21] ),
    .X(\CPU_imem_rd_data_a1[23] ));
 sky130_fd_sc_hd__o31ai_1 _10119_ (.A1(_01148_),
    .A2(_01151_),
    .A3(_04223_),
    .B1(_04222_),
    .Y(\CPU_imm_a1[3] ));
 sky130_fd_sc_hd__a21boi_1 _10120_ (.A1(_01156_),
    .A2(_01149_),
    .B1_N(net1833),
    .Y(_04224_));
 sky130_fd_sc_hd__nor3_1 _10121_ (.A(\CPU_dec_bits_a1[10] ),
    .B(_01148_),
    .C(_04224_),
    .Y(CPU_is_add_a1));
 sky130_fd_sc_hd__nor3b_1 _10122_ (.A(\CPU_imm_a1[10] ),
    .B(_04224_),
    .C_N(_01148_),
    .Y(CPU_is_addi_a1));
 sky130_fd_sc_hd__nor4_1 _10123_ (.A(_05822_),
    .B(_05817_),
    .C(_05820_),
    .D(_01122_),
    .Y(CPU_is_blt_a1));
 sky130_fd_sc_hd__nor2_1 _10124_ (.A(\CPU_dec_bits_a1[10] ),
    .B(_01152_),
    .Y(CPU_rd_valid_a1));
 sky130_fd_sc_hd__inv_1 _10125_ (.A(_03217_),
    .Y(\CPU_result_a3[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_163 ();
 sky130_fd_sc_hd__nor2_2 _10128_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .Y(_04227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_161 ();
 sky130_fd_sc_hd__nor2_2 _10131_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_8 _10132_ (.A(_04227_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_160 ();
 sky130_fd_sc_hd__nand2_8 _10134_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04233_));
 sky130_fd_sc_hd__nor3_4 _10135_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .C(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__nor4_4 _10138_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .C(\CPU_rf_rd_index1_a2[1] ),
    .D(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__a21oi_1 _10140_ (.A1(\CPU_Xreg_value_a4[3][0] ),
    .A2(net40),
    .B1(net93),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2b_4 _10141_ (.A_N(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04240_));
 sky130_fd_sc_hd__nor3_4 _10142_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .C(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__nand2b_4 _10145_ (.A_N(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .Y(_04244_));
 sky130_fd_sc_hd__nor3_4 _10146_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .C(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_153 ();
 sky130_fd_sc_hd__a22oi_1 _10149_ (.A1(\CPU_Xreg_value_a4[1][0] ),
    .A2(net37),
    .B1(_04245_),
    .B2(\CPU_Xreg_value_a4[8][0] ),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_8 _10150_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .Y(_04249_));
 sky130_fd_sc_hd__nor2_8 _10151_ (.A(_04240_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_152 ();
 sky130_fd_sc_hd__nor2_8 _10153_ (.A(_04240_),
    .B(_04244_),
    .Y(_04252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__a22oi_1 _10156_ (.A1(\CPU_Xreg_value_a4[13][0] ),
    .A2(_04250_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][0] ),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2b_4 _10157_ (.A_N(\CPU_rf_rd_index1_a2[3] ),
    .B(\CPU_rf_rd_index1_a2[2] ),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2b_4 _10158_ (.A_N(\CPU_rf_rd_index1_a2[0] ),
    .B(\CPU_rf_rd_index1_a2[1] ),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_8 _10159_ (.A(_04256_),
    .B(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__nor2_8 _10161_ (.A(_04256_),
    .B(_04233_),
    .Y(_04260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_148 ();
 sky130_fd_sc_hd__a22oi_1 _10163_ (.A1(\CPU_Xreg_value_a4[6][0] ),
    .A2(_04258_),
    .B1(_04260_),
    .B2(\CPU_Xreg_value_a4[7][0] ),
    .Y(_04262_));
 sky130_fd_sc_hd__nand4_1 _10164_ (.A(_04239_),
    .B(_04248_),
    .C(_04255_),
    .D(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__nor3_4 _10165_ (.A(\CPU_rf_rd_index1_a2[2] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .C(_04257_),
    .Y(_04264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_147 ();
 sky130_fd_sc_hd__nor3_4 _10167_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .C(_04249_),
    .Y(_04266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_146 ();
 sky130_fd_sc_hd__nor2_8 _10169_ (.A(_04233_),
    .B(_04249_),
    .Y(_04268_));
 sky130_fd_sc_hd__nor3_4 _10170_ (.A(\CPU_rf_rd_index1_a2[1] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .C(_04256_),
    .Y(_04269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_145 ();
 sky130_fd_sc_hd__a22o_1 _10172_ (.A1(\CPU_Xreg_value_a4[15][0] ),
    .A2(_04268_),
    .B1(net28),
    .B2(\CPU_Xreg_value_a4[4][0] ),
    .X(_04271_));
 sky130_fd_sc_hd__a221oi_1 _10173_ (.A1(\CPU_Xreg_value_a4[2][0] ),
    .A2(_04264_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][0] ),
    .C1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__nor2_8 _10174_ (.A(_04257_),
    .B(_04244_),
    .Y(_04273_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_144 ();
 sky130_fd_sc_hd__nor2_8 _10176_ (.A(_04233_),
    .B(_04244_),
    .Y(_04275_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__a22oi_1 _10179_ (.A1(\CPU_Xreg_value_a4[10][0] ),
    .A2(_04273_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][0] ),
    .Y(_04278_));
 sky130_fd_sc_hd__nor2_8 _10180_ (.A(_04257_),
    .B(_04249_),
    .Y(_04279_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__nor2_8 _10182_ (.A(_04240_),
    .B(_04256_),
    .Y(_04281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_140 ();
 sky130_fd_sc_hd__a22oi_1 _10184_ (.A1(\CPU_Xreg_value_a4[14][0] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][0] ),
    .Y(_04283_));
 sky130_fd_sc_hd__nand3_1 _10185_ (.A(_04272_),
    .B(_04278_),
    .C(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__o22ai_4 _10186_ (.A1(\CPU_Xreg_value_a4[0][0] ),
    .A2(_04231_),
    .B1(_04263_),
    .B2(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21o_2 _10187_ (.A1(_02568_),
    .A2(_02573_),
    .B1(\CPU_rd_a3[4] ),
    .X(_04286_));
 sky130_fd_sc_hd__xnor2_1 _10188_ (.A(\CPU_rd_a3[3] ),
    .B(\CPU_rf_rd_index1_a2[3] ),
    .Y(_04287_));
 sky130_fd_sc_hd__xnor2_1 _10189_ (.A(\CPU_rd_a3[2] ),
    .B(\CPU_rf_rd_index1_a2[2] ),
    .Y(_04288_));
 sky130_fd_sc_hd__xnor2_1 _10190_ (.A(\CPU_rd_a3[0] ),
    .B(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04289_));
 sky130_fd_sc_hd__xnor2_1 _10191_ (.A(\CPU_rd_a3[1] ),
    .B(\CPU_rf_rd_index1_a2[1] ),
    .Y(_04290_));
 sky130_fd_sc_hd__nand4_4 _10192_ (.A(_04287_),
    .B(_04288_),
    .C(_04289_),
    .D(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__nor2_8 _10193_ (.A(_04286_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_139 ();
 sky130_fd_sc_hd__mux2i_4 _10195_ (.A0(_04285_),
    .A1(_02560_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[0] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 ();
 sky130_fd_sc_hd__a21oi_1 _10199_ (.A1(net1236),
    .A2(net31),
    .B1(net94),
    .Y(_04297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_134 ();
 sky130_fd_sc_hd__a22oi_1 _10202_ (.A1(\CPU_Xreg_value_a4[14][10] ),
    .A2(_04279_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][10] ),
    .Y(_04300_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_132 ();
 sky130_fd_sc_hd__a22oi_1 _10205_ (.A1(\CPU_Xreg_value_a4[13][10] ),
    .A2(_04250_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][10] ),
    .Y(_04303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_130 ();
 sky130_fd_sc_hd__a22oi_1 _10208_ (.A1(\CPU_Xreg_value_a4[6][10] ),
    .A2(_04258_),
    .B1(net29),
    .B2(net1347),
    .Y(_04306_));
 sky130_fd_sc_hd__nand4_1 _10209_ (.A(_04297_),
    .B(_04300_),
    .C(_04303_),
    .D(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_128 ();
 sky130_fd_sc_hd__a22o_1 _10212_ (.A1(\CPU_Xreg_value_a4[11][10] ),
    .A2(_04275_),
    .B1(net40),
    .B2(\CPU_Xreg_value_a4[3][10] ),
    .X(_04310_));
 sky130_fd_sc_hd__a221oi_1 _10213_ (.A1(net1253),
    .A2(_04260_),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][10] ),
    .C1(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__a22oi_1 _10216_ (.A1(\CPU_Xreg_value_a4[1][10] ),
    .A2(net36),
    .B1(net33),
    .B2(\CPU_Xreg_value_a4[2][10] ),
    .Y(_04314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__a22oi_1 _10220_ (.A1(net1717),
    .A2(net34),
    .B1(_04268_),
    .B2(net1278),
    .Y(_04318_));
 sky130_fd_sc_hd__nand3_1 _10221_ (.A(_04311_),
    .B(_04314_),
    .C(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__o22ai_1 _10222_ (.A1(net1292),
    .A2(_04231_),
    .B1(_04307_),
    .B2(net1718),
    .Y(_04320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__nand2_1 _10224_ (.A(_02635_),
    .B(_04292_),
    .Y(_04322_));
 sky130_fd_sc_hd__o21ai_0 _10225_ (.A1(_04292_),
    .A2(_04320_),
    .B1(_04322_),
    .Y(\CPU_src1_value_a2[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_121 ();
 sky130_fd_sc_hd__a21oi_1 _10227_ (.A1(\CPU_Xreg_value_a4[4][11] ),
    .A2(net27),
    .B1(net93),
    .Y(_04324_));
 sky130_fd_sc_hd__a22oi_1 _10228_ (.A1(\CPU_Xreg_value_a4[6][11] ),
    .A2(_04258_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][11] ),
    .Y(_04325_));
 sky130_fd_sc_hd__a22oi_1 _10229_ (.A1(\CPU_Xreg_value_a4[10][11] ),
    .A2(_04273_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][11] ),
    .Y(_04326_));
 sky130_fd_sc_hd__a22oi_1 _10230_ (.A1(\CPU_Xreg_value_a4[11][11] ),
    .A2(_04275_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][11] ),
    .Y(_04327_));
 sky130_fd_sc_hd__nand4_2 _10231_ (.A(_04324_),
    .B(_04325_),
    .C(_04326_),
    .D(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__a22o_1 _10232_ (.A1(\CPU_Xreg_value_a4[7][11] ),
    .A2(_04260_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][11] ),
    .X(_04329_));
 sky130_fd_sc_hd__a221oi_1 _10233_ (.A1(\CPU_Xreg_value_a4[1][11] ),
    .A2(net36),
    .B1(net34),
    .B2(\CPU_Xreg_value_a4[8][11] ),
    .C1(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__a22oi_1 _10236_ (.A1(\CPU_Xreg_value_a4[2][11] ),
    .A2(net32),
    .B1(net31),
    .B2(\CPU_Xreg_value_a4[12][11] ),
    .Y(_04333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__a22oi_1 _10238_ (.A1(\CPU_Xreg_value_a4[14][11] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][11] ),
    .Y(_04335_));
 sky130_fd_sc_hd__nand3_1 _10239_ (.A(_04330_),
    .B(_04333_),
    .C(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__o22ai_4 _10240_ (.A1(net1504),
    .A2(_04231_),
    .B1(_04328_),
    .B2(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand3_1 _10241_ (.A(_02661_),
    .B(_02678_),
    .C(_02681_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(_04338_),
    .B(_04292_),
    .Y(_04339_));
 sky130_fd_sc_hd__o21ai_0 _10243_ (.A1(_04292_),
    .A2(_04337_),
    .B1(_04339_),
    .Y(\CPU_src1_value_a2[11] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__a21oi_1 _10245_ (.A1(\CPU_Xreg_value_a4[3][12] ),
    .A2(_04234_),
    .B1(net95),
    .Y(_04341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__a22oi_1 _10247_ (.A1(\CPU_Xreg_value_a4[1][12] ),
    .A2(_04241_),
    .B1(_04245_),
    .B2(\CPU_Xreg_value_a4[8][12] ),
    .Y(_04343_));
 sky130_fd_sc_hd__a22oi_1 _10248_ (.A1(\CPU_Xreg_value_a4[13][12] ),
    .A2(_04250_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][12] ),
    .Y(_04344_));
 sky130_fd_sc_hd__a22oi_1 _10249_ (.A1(\CPU_Xreg_value_a4[14][12] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][12] ),
    .Y(_04345_));
 sky130_fd_sc_hd__nand4_1 _10250_ (.A(_04341_),
    .B(_04343_),
    .C(_04344_),
    .D(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__a22o_1 _10251_ (.A1(\CPU_Xreg_value_a4[12][12] ),
    .A2(_04266_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][12] ),
    .X(_04347_));
 sky130_fd_sc_hd__a221oi_1 _10252_ (.A1(\CPU_Xreg_value_a4[6][12] ),
    .A2(_04258_),
    .B1(_04264_),
    .B2(\CPU_Xreg_value_a4[2][12] ),
    .C1(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_115 ();
 sky130_fd_sc_hd__a22oi_1 _10254_ (.A1(\CPU_Xreg_value_a4[7][12] ),
    .A2(_04260_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][12] ),
    .Y(_04350_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_114 ();
 sky130_fd_sc_hd__a22oi_1 _10256_ (.A1(\CPU_Xreg_value_a4[10][12] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][12] ),
    .Y(_04352_));
 sky130_fd_sc_hd__nand3_1 _10257_ (.A(_04348_),
    .B(_04350_),
    .C(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__o22ai_4 _10258_ (.A1(\CPU_Xreg_value_a4[0][12] ),
    .A2(_04231_),
    .B1(_04346_),
    .B2(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand2_1 _10259_ (.A(_02710_),
    .B(_04292_),
    .Y(_04355_));
 sky130_fd_sc_hd__o21ai_0 _10260_ (.A1(_04292_),
    .A2(_04354_),
    .B1(_04355_),
    .Y(\CPU_src1_value_a2[12] ));
 sky130_fd_sc_hd__a21oi_1 _10261_ (.A1(\CPU_Xreg_value_a4[12][13] ),
    .A2(net31),
    .B1(net94),
    .Y(_04356_));
 sky130_fd_sc_hd__a22oi_1 _10262_ (.A1(\CPU_Xreg_value_a4[1][13] ),
    .A2(net36),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][13] ),
    .Y(_04357_));
 sky130_fd_sc_hd__a22oi_1 _10263_ (.A1(\CPU_Xreg_value_a4[13][13] ),
    .A2(_04250_),
    .B1(net38),
    .B2(\CPU_Xreg_value_a4[3][13] ),
    .Y(_04358_));
 sky130_fd_sc_hd__a22oi_1 _10264_ (.A1(\CPU_Xreg_value_a4[14][13] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][13] ),
    .Y(_04359_));
 sky130_fd_sc_hd__nand4_2 _10265_ (.A(_04356_),
    .B(_04357_),
    .C(_04358_),
    .D(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_113 ();
 sky130_fd_sc_hd__a22oi_1 _10267_ (.A1(\CPU_Xreg_value_a4[6][13] ),
    .A2(_04258_),
    .B1(net33),
    .B2(\CPU_Xreg_value_a4[2][13] ),
    .Y(_04362_));
 sky130_fd_sc_hd__a22oi_1 _10268_ (.A1(\CPU_Xreg_value_a4[4][13] ),
    .A2(net28),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][13] ),
    .Y(_04363_));
 sky130_fd_sc_hd__a22oi_1 _10269_ (.A1(\CPU_Xreg_value_a4[7][13] ),
    .A2(_04260_),
    .B1(net34),
    .B2(\CPU_Xreg_value_a4[8][13] ),
    .Y(_04364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_112 ();
 sky130_fd_sc_hd__a22oi_1 _10271_ (.A1(\CPU_Xreg_value_a4[10][13] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][13] ),
    .Y(_04366_));
 sky130_fd_sc_hd__nand4_1 _10272_ (.A(_04362_),
    .B(_04363_),
    .C(_04364_),
    .D(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__o22ai_4 _10273_ (.A1(\CPU_Xreg_value_a4[0][13] ),
    .A2(_04231_),
    .B1(_04360_),
    .B2(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__and2_1 _10274_ (.A(_02735_),
    .B(_02746_),
    .X(_04369_));
 sky130_fd_sc_hd__mux2i_4 _10275_ (.A0(_04368_),
    .A1(_04369_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[13] ));
 sky130_fd_sc_hd__a21oi_1 _10276_ (.A1(net1744),
    .A2(net31),
    .B1(_04237_),
    .Y(_04370_));
 sky130_fd_sc_hd__a22oi_1 _10277_ (.A1(\CPU_Xreg_value_a4[2][14] ),
    .A2(net33),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][14] ),
    .Y(_04371_));
 sky130_fd_sc_hd__a22oi_1 _10278_ (.A1(\CPU_Xreg_value_a4[6][14] ),
    .A2(_04258_),
    .B1(net40),
    .B2(\CPU_Xreg_value_a4[3][14] ),
    .Y(_04372_));
 sky130_fd_sc_hd__a22oi_1 _10279_ (.A1(\CPU_Xreg_value_a4[10][14] ),
    .A2(_04273_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][14] ),
    .Y(_04373_));
 sky130_fd_sc_hd__nand4_1 _10280_ (.A(_04370_),
    .B(_04371_),
    .C(_04372_),
    .D(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a22oi_1 _10281_ (.A1(\CPU_Xreg_value_a4[7][14] ),
    .A2(_04260_),
    .B1(_04252_),
    .B2(net1365),
    .Y(_04375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_111 ();
 sky130_fd_sc_hd__a22oi_1 _10283_ (.A1(\CPU_Xreg_value_a4[14][14] ),
    .A2(_04279_),
    .B1(net29),
    .B2(\CPU_Xreg_value_a4[4][14] ),
    .Y(_04377_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_110 ();
 sky130_fd_sc_hd__a22oi_1 _10285_ (.A1(\CPU_Xreg_value_a4[1][14] ),
    .A2(net37),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][14] ),
    .Y(_04379_));
 sky130_fd_sc_hd__a22oi_1 _10286_ (.A1(\CPU_Xreg_value_a4[8][14] ),
    .A2(_04245_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][14] ),
    .Y(_04380_));
 sky130_fd_sc_hd__nand4_1 _10287_ (.A(_04375_),
    .B(_04377_),
    .C(_04379_),
    .D(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__o22ai_1 _10288_ (.A1(net1269),
    .A2(_04231_),
    .B1(net1745),
    .B2(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__mux2i_1 _10289_ (.A0(_04382_),
    .A1(_02764_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[14] ));
 sky130_fd_sc_hd__a22o_1 _10290_ (.A1(\CPU_Xreg_value_a4[6][15] ),
    .A2(_04258_),
    .B1(net31),
    .B2(\CPU_Xreg_value_a4[12][15] ),
    .X(_04383_));
 sky130_fd_sc_hd__a221oi_1 _10291_ (.A1(\CPU_Xreg_value_a4[7][15] ),
    .A2(_04260_),
    .B1(net29),
    .B2(\CPU_Xreg_value_a4[4][15] ),
    .C1(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a22o_1 _10292_ (.A1(\CPU_Xreg_value_a4[8][15] ),
    .A2(_04245_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][15] ),
    .X(_04385_));
 sky130_fd_sc_hd__a221oi_1 _10293_ (.A1(\CPU_Xreg_value_a4[10][15] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][15] ),
    .C1(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__mux2i_1 _10294_ (.A0(\CPU_Xreg_value_a4[2][15] ),
    .A1(\CPU_Xreg_value_a4[3][15] ),
    .S(\CPU_rf_rd_index1_a2[0] ),
    .Y(_04387_));
 sky130_fd_sc_hd__o21ai_0 _10295_ (.A1(\CPU_Xreg_value_a4[1][15] ),
    .A2(_04240_),
    .B1(_04227_),
    .Y(_04388_));
 sky130_fd_sc_hd__a21oi_1 _10296_ (.A1(\CPU_rf_rd_index1_a2[1] ),
    .A2(_04387_),
    .B1(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__a221o_1 _10297_ (.A1(\CPU_Xreg_value_a4[13][15] ),
    .A2(_04250_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][15] ),
    .C1(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__a221oi_2 _10298_ (.A1(\CPU_Xreg_value_a4[11][15] ),
    .A2(_04275_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][15] ),
    .C1(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand3_1 _10299_ (.A(_04384_),
    .B(_04386_),
    .C(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__o21ai_1 _10300_ (.A1(net1307),
    .A2(_04231_),
    .B1(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_02782_),
    .B(_04292_),
    .Y(_04394_));
 sky130_fd_sc_hd__o21ai_0 _10302_ (.A1(_04292_),
    .A2(_04393_),
    .B1(_04394_),
    .Y(\CPU_src1_value_a2[15] ));
 sky130_fd_sc_hd__a21oi_1 _10303_ (.A1(\CPU_Xreg_value_a4[4][16] ),
    .A2(net29),
    .B1(_04237_),
    .Y(_04395_));
 sky130_fd_sc_hd__a22oi_1 _10304_ (.A1(\CPU_Xreg_value_a4[2][16] ),
    .A2(net33),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][16] ),
    .Y(_04396_));
 sky130_fd_sc_hd__a22oi_1 _10305_ (.A1(\CPU_Xreg_value_a4[8][16] ),
    .A2(_04245_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][16] ),
    .Y(_04397_));
 sky130_fd_sc_hd__a22oi_1 _10306_ (.A1(\CPU_Xreg_value_a4[10][16] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][16] ),
    .Y(_04398_));
 sky130_fd_sc_hd__nand4_1 _10307_ (.A(_04395_),
    .B(_04396_),
    .C(_04397_),
    .D(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__a22oi_1 _10308_ (.A1(\CPU_Xreg_value_a4[1][16] ),
    .A2(net37),
    .B1(net31),
    .B2(\CPU_Xreg_value_a4[12][16] ),
    .Y(_04400_));
 sky130_fd_sc_hd__a22oi_1 _10309_ (.A1(\CPU_Xreg_value_a4[13][16] ),
    .A2(_04250_),
    .B1(net40),
    .B2(net1797),
    .Y(_04401_));
 sky130_fd_sc_hd__a22oi_1 _10310_ (.A1(\CPU_Xreg_value_a4[6][16] ),
    .A2(_04258_),
    .B1(_04260_),
    .B2(\CPU_Xreg_value_a4[7][16] ),
    .Y(_04402_));
 sky130_fd_sc_hd__a22oi_1 _10311_ (.A1(\CPU_Xreg_value_a4[14][16] ),
    .A2(_04279_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][16] ),
    .Y(_04403_));
 sky130_fd_sc_hd__nand4_1 _10312_ (.A(_04400_),
    .B(_04401_),
    .C(_04402_),
    .D(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__o22ai_1 _10313_ (.A1(net1312),
    .A2(_04231_),
    .B1(_04399_),
    .B2(net1798),
    .Y(_04405_));
 sky130_fd_sc_hd__mux2i_1 _10314_ (.A0(net1799),
    .A1(_02807_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[16] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_109 ();
 sky130_fd_sc_hd__a21oi_1 _10316_ (.A1(\CPU_Xreg_value_a4[14][17] ),
    .A2(_04279_),
    .B1(net93),
    .Y(_04407_));
 sky130_fd_sc_hd__a22oi_1 _10317_ (.A1(\CPU_Xreg_value_a4[10][17] ),
    .A2(_04273_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][17] ),
    .Y(_04408_));
 sky130_fd_sc_hd__a22oi_1 _10318_ (.A1(\CPU_Xreg_value_a4[2][17] ),
    .A2(_04264_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][17] ),
    .Y(_04409_));
 sky130_fd_sc_hd__a22oi_1 _10319_ (.A1(\CPU_Xreg_value_a4[4][17] ),
    .A2(net28),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][17] ),
    .Y(_04410_));
 sky130_fd_sc_hd__nand4_1 _10320_ (.A(_04407_),
    .B(_04408_),
    .C(_04409_),
    .D(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__a22o_1 _10321_ (.A1(\CPU_Xreg_value_a4[1][17] ),
    .A2(net37),
    .B1(net38),
    .B2(\CPU_Xreg_value_a4[3][17] ),
    .X(_04412_));
 sky130_fd_sc_hd__a221oi_1 _10322_ (.A1(\CPU_Xreg_value_a4[6][17] ),
    .A2(_04258_),
    .B1(_04245_),
    .B2(\CPU_Xreg_value_a4[8][17] ),
    .C1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_108 ();
 sky130_fd_sc_hd__a22oi_1 _10324_ (.A1(\CPU_Xreg_value_a4[11][17] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][17] ),
    .Y(_04415_));
 sky130_fd_sc_hd__a22oi_1 _10325_ (.A1(\CPU_Xreg_value_a4[7][17] ),
    .A2(_04260_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][17] ),
    .Y(_04416_));
 sky130_fd_sc_hd__nand3_1 _10326_ (.A(_04413_),
    .B(_04415_),
    .C(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__o22ai_2 _10327_ (.A1(net1418),
    .A2(_04231_),
    .B1(_04411_),
    .B2(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_107 ();
 sky130_fd_sc_hd__mux2i_1 _10329_ (.A0(_04418_),
    .A1(_02832_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[17] ));
 sky130_fd_sc_hd__a22oi_1 _10330_ (.A1(\CPU_Xreg_value_a4[13][18] ),
    .A2(_04250_),
    .B1(net40),
    .B2(\CPU_Xreg_value_a4[3][18] ),
    .Y(_04420_));
 sky130_fd_sc_hd__a22oi_1 _10331_ (.A1(\CPU_Xreg_value_a4[10][18] ),
    .A2(_04273_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][18] ),
    .Y(_04421_));
 sky130_fd_sc_hd__a22oi_1 _10332_ (.A1(\CPU_Xreg_value_a4[8][18] ),
    .A2(net34),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][18] ),
    .Y(_04422_));
 sky130_fd_sc_hd__a22oi_1 _10333_ (.A1(\CPU_Xreg_value_a4[6][18] ),
    .A2(_04258_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][18] ),
    .Y(_04423_));
 sky130_fd_sc_hd__nand4_1 _10334_ (.A(_04420_),
    .B(_04421_),
    .C(_04422_),
    .D(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__a22oi_1 _10335_ (.A1(\CPU_Xreg_value_a4[7][18] ),
    .A2(_04260_),
    .B1(net29),
    .B2(net1845),
    .Y(_04425_));
 sky130_fd_sc_hd__a22oi_1 _10336_ (.A1(\CPU_Xreg_value_a4[1][18] ),
    .A2(net36),
    .B1(net31),
    .B2(net1710),
    .Y(_04426_));
 sky130_fd_sc_hd__a22oi_1 _10337_ (.A1(\CPU_Xreg_value_a4[2][18] ),
    .A2(net33),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][18] ),
    .Y(_04427_));
 sky130_fd_sc_hd__a21oi_1 _10338_ (.A1(\CPU_Xreg_value_a4[14][18] ),
    .A2(_04279_),
    .B1(net94),
    .Y(_04428_));
 sky130_fd_sc_hd__nand4_1 _10339_ (.A(net1846),
    .B(_04426_),
    .C(_04427_),
    .D(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__o22ai_2 _10340_ (.A1(net1610),
    .A2(_04231_),
    .B1(_04424_),
    .B2(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__mux2i_1 _10341_ (.A0(_04430_),
    .A1(_02853_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[18] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_106 ();
 sky130_fd_sc_hd__a21oi_1 _10343_ (.A1(\CPU_Xreg_value_a4[2][19] ),
    .A2(_04264_),
    .B1(net93),
    .Y(_04432_));
 sky130_fd_sc_hd__a22oi_1 _10344_ (.A1(\CPU_Xreg_value_a4[1][19] ),
    .A2(net37),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][19] ),
    .Y(_04433_));
 sky130_fd_sc_hd__a22oi_1 _10345_ (.A1(\CPU_Xreg_value_a4[10][19] ),
    .A2(_04273_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][19] ),
    .Y(_04434_));
 sky130_fd_sc_hd__a22oi_1 _10346_ (.A1(\CPU_Xreg_value_a4[12][19] ),
    .A2(net30),
    .B1(net28),
    .B2(\CPU_Xreg_value_a4[4][19] ),
    .Y(_04435_));
 sky130_fd_sc_hd__nand4_1 _10347_ (.A(_04432_),
    .B(_04433_),
    .C(_04434_),
    .D(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__a22o_1 _10348_ (.A1(\CPU_Xreg_value_a4[3][19] ),
    .A2(net38),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][19] ),
    .X(_04437_));
 sky130_fd_sc_hd__a221oi_1 _10349_ (.A1(net1750),
    .A2(_04260_),
    .B1(_04245_),
    .B2(net1735),
    .C1(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__a22oi_1 _10350_ (.A1(\CPU_Xreg_value_a4[6][19] ),
    .A2(_04258_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][19] ),
    .Y(_04439_));
 sky130_fd_sc_hd__a22oi_1 _10351_ (.A1(\CPU_Xreg_value_a4[13][19] ),
    .A2(_04250_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][19] ),
    .Y(_04440_));
 sky130_fd_sc_hd__nand3_1 _10352_ (.A(_04438_),
    .B(_04439_),
    .C(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o22ai_2 _10353_ (.A1(net1409),
    .A2(_04231_),
    .B1(_04436_),
    .B2(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__o21ai_0 _10354_ (.A1(_02866_),
    .A2(_02881_),
    .B1(_04292_),
    .Y(_04443_));
 sky130_fd_sc_hd__o21ai_0 _10355_ (.A1(_04292_),
    .A2(_04442_),
    .B1(_04443_),
    .Y(\CPU_src1_value_a2[19] ));
 sky130_fd_sc_hd__a21oi_1 _10356_ (.A1(\CPU_Xreg_value_a4[2][1] ),
    .A2(_04264_),
    .B1(net95),
    .Y(_04444_));
 sky130_fd_sc_hd__a22oi_1 _10357_ (.A1(\CPU_Xreg_value_a4[12][1] ),
    .A2(_04266_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][1] ),
    .Y(_04445_));
 sky130_fd_sc_hd__a22oi_1 _10358_ (.A1(\CPU_Xreg_value_a4[6][1] ),
    .A2(_04258_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][1] ),
    .Y(_04446_));
 sky130_fd_sc_hd__a22oi_1 _10359_ (.A1(\CPU_Xreg_value_a4[3][1] ),
    .A2(_04234_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][1] ),
    .Y(_04447_));
 sky130_fd_sc_hd__nand4_2 _10360_ (.A(_04444_),
    .B(_04445_),
    .C(_04446_),
    .D(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__a22o_1 _10361_ (.A1(\CPU_Xreg_value_a4[1][1] ),
    .A2(_04241_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][1] ),
    .X(_04449_));
 sky130_fd_sc_hd__a221oi_1 _10362_ (.A1(\CPU_Xreg_value_a4[11][1] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][1] ),
    .C1(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__a22oi_1 _10363_ (.A1(\CPU_Xreg_value_a4[10][1] ),
    .A2(_04273_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][1] ),
    .Y(_04451_));
 sky130_fd_sc_hd__a22oi_1 _10364_ (.A1(\CPU_Xreg_value_a4[7][1] ),
    .A2(_04260_),
    .B1(net35),
    .B2(\CPU_Xreg_value_a4[8][1] ),
    .Y(_04452_));
 sky130_fd_sc_hd__nand3_1 _10365_ (.A(_04450_),
    .B(_04451_),
    .C(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__o22ai_4 _10366_ (.A1(net1855),
    .A2(_04231_),
    .B1(_04448_),
    .B2(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _10367_ (.A(_02888_),
    .B(_04292_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ai_0 _10368_ (.A1(_04292_),
    .A2(_04454_),
    .B1(_04455_),
    .Y(\CPU_src1_value_a2[1] ));
 sky130_fd_sc_hd__a21oi_1 _10369_ (.A1(\CPU_Xreg_value_a4[2][20] ),
    .A2(_04264_),
    .B1(net93),
    .Y(_04456_));
 sky130_fd_sc_hd__a22oi_1 _10370_ (.A1(\CPU_Xreg_value_a4[7][20] ),
    .A2(_04260_),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][20] ),
    .Y(_04457_));
 sky130_fd_sc_hd__a22oi_1 _10371_ (.A1(\CPU_Xreg_value_a4[13][20] ),
    .A2(_04250_),
    .B1(net27),
    .B2(\CPU_Xreg_value_a4[4][20] ),
    .Y(_04458_));
 sky130_fd_sc_hd__a22oi_1 _10372_ (.A1(\CPU_Xreg_value_a4[12][20] ),
    .A2(net30),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][20] ),
    .Y(_04459_));
 sky130_fd_sc_hd__nand4_2 _10373_ (.A(_04456_),
    .B(_04457_),
    .C(_04458_),
    .D(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__a22o_1 _10374_ (.A1(\CPU_Xreg_value_a4[8][20] ),
    .A2(net35),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][20] ),
    .X(_04461_));
 sky130_fd_sc_hd__a221oi_1 _10375_ (.A1(\CPU_Xreg_value_a4[1][20] ),
    .A2(net37),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][20] ),
    .C1(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__a22oi_1 _10376_ (.A1(\CPU_Xreg_value_a4[6][20] ),
    .A2(_04258_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][20] ),
    .Y(_04463_));
 sky130_fd_sc_hd__a22oi_1 _10377_ (.A1(\CPU_Xreg_value_a4[15][20] ),
    .A2(_04268_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][20] ),
    .Y(_04464_));
 sky130_fd_sc_hd__nand3_1 _10378_ (.A(_04462_),
    .B(_04463_),
    .C(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__o22ai_4 _10379_ (.A1(net1675),
    .A2(_04231_),
    .B1(_04460_),
    .B2(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__mux2i_1 _10380_ (.A0(_04466_),
    .A1(_02908_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[20] ));
 sky130_fd_sc_hd__a21oi_1 _10381_ (.A1(\CPU_Xreg_value_a4[11][21] ),
    .A2(_04275_),
    .B1(net95),
    .Y(_04467_));
 sky130_fd_sc_hd__a22oi_1 _10382_ (.A1(\CPU_Xreg_value_a4[4][21] ),
    .A2(net27),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][21] ),
    .Y(_04468_));
 sky130_fd_sc_hd__a22oi_1 _10383_ (.A1(\CPU_Xreg_value_a4[10][21] ),
    .A2(_04273_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][21] ),
    .Y(_04469_));
 sky130_fd_sc_hd__a22oi_1 _10384_ (.A1(\CPU_Xreg_value_a4[1][21] ),
    .A2(net37),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][21] ),
    .Y(_04470_));
 sky130_fd_sc_hd__nand4_1 _10385_ (.A(_04467_),
    .B(_04468_),
    .C(_04469_),
    .D(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__a22o_1 _10386_ (.A1(\CPU_Xreg_value_a4[2][21] ),
    .A2(net32),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][21] ),
    .X(_04472_));
 sky130_fd_sc_hd__a221oi_1 _10387_ (.A1(\CPU_Xreg_value_a4[7][21] ),
    .A2(_04260_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][21] ),
    .C1(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a22oi_1 _10388_ (.A1(\CPU_Xreg_value_a4[6][21] ),
    .A2(_04258_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][21] ),
    .Y(_04474_));
 sky130_fd_sc_hd__a22oi_1 _10389_ (.A1(\CPU_Xreg_value_a4[8][21] ),
    .A2(net35),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][21] ),
    .Y(_04475_));
 sky130_fd_sc_hd__nand3_1 _10390_ (.A(_04473_),
    .B(_04474_),
    .C(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__o22ai_4 _10391_ (.A1(net1671),
    .A2(_04231_),
    .B1(_04471_),
    .B2(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__mux2i_1 _10392_ (.A0(_04477_),
    .A1(_02934_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[21] ));
 sky130_fd_sc_hd__a21oi_1 _10393_ (.A1(\CPU_Xreg_value_a4[12][22] ),
    .A2(net31),
    .B1(net94),
    .Y(_04478_));
 sky130_fd_sc_hd__a22oi_1 _10394_ (.A1(\CPU_Xreg_value_a4[11][22] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][22] ),
    .Y(_04479_));
 sky130_fd_sc_hd__a22oi_1 _10395_ (.A1(\CPU_Xreg_value_a4[10][22] ),
    .A2(_04273_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][22] ),
    .Y(_04480_));
 sky130_fd_sc_hd__a22oi_1 _10396_ (.A1(\CPU_Xreg_value_a4[4][22] ),
    .A2(net28),
    .B1(net38),
    .B2(\CPU_Xreg_value_a4[3][22] ),
    .Y(_04481_));
 sky130_fd_sc_hd__nand4_1 _10397_ (.A(_04478_),
    .B(_04479_),
    .C(_04480_),
    .D(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__a22o_1 _10398_ (.A1(\CPU_Xreg_value_a4[2][22] ),
    .A2(net33),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][22] ),
    .X(_04483_));
 sky130_fd_sc_hd__a221oi_1 _10399_ (.A1(\CPU_Xreg_value_a4[1][22] ),
    .A2(net36),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][22] ),
    .C1(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a22oi_1 _10400_ (.A1(\CPU_Xreg_value_a4[8][22] ),
    .A2(net34),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][22] ),
    .Y(_04485_));
 sky130_fd_sc_hd__a22oi_1 _10401_ (.A1(\CPU_Xreg_value_a4[6][22] ),
    .A2(_04258_),
    .B1(_04260_),
    .B2(\CPU_Xreg_value_a4[7][22] ),
    .Y(_04486_));
 sky130_fd_sc_hd__nand3_1 _10402_ (.A(_04484_),
    .B(_04485_),
    .C(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__o22ai_2 _10403_ (.A1(net1607),
    .A2(_04231_),
    .B1(_04482_),
    .B2(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__mux2i_1 _10404_ (.A0(_04488_),
    .A1(_02959_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[22] ));
 sky130_fd_sc_hd__a21oi_1 _10405_ (.A1(\CPU_Xreg_value_a4[15][23] ),
    .A2(_04268_),
    .B1(net93),
    .Y(_04489_));
 sky130_fd_sc_hd__a22oi_1 _10406_ (.A1(\CPU_Xreg_value_a4[7][23] ),
    .A2(_04260_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][23] ),
    .Y(_04490_));
 sky130_fd_sc_hd__a22oi_1 _10407_ (.A1(\CPU_Xreg_value_a4[8][23] ),
    .A2(net35),
    .B1(net27),
    .B2(\CPU_Xreg_value_a4[4][23] ),
    .Y(_04491_));
 sky130_fd_sc_hd__a22oi_1 _10408_ (.A1(\CPU_Xreg_value_a4[11][23] ),
    .A2(_04275_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][23] ),
    .Y(_04492_));
 sky130_fd_sc_hd__nand4_1 _10409_ (.A(_04489_),
    .B(_04490_),
    .C(_04491_),
    .D(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__a22o_1 _10410_ (.A1(\CPU_Xreg_value_a4[2][23] ),
    .A2(net32),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][23] ),
    .X(_04494_));
 sky130_fd_sc_hd__a221oi_1 _10411_ (.A1(\CPU_Xreg_value_a4[1][23] ),
    .A2(net37),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][23] ),
    .C1(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__a22oi_1 _10412_ (.A1(\CPU_Xreg_value_a4[10][23] ),
    .A2(_04273_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][23] ),
    .Y(_04496_));
 sky130_fd_sc_hd__a22oi_1 _10413_ (.A1(\CPU_Xreg_value_a4[6][23] ),
    .A2(_04258_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][23] ),
    .Y(_04497_));
 sky130_fd_sc_hd__nand3_1 _10414_ (.A(_04495_),
    .B(_04496_),
    .C(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__o22ai_4 _10415_ (.A1(net1511),
    .A2(_04231_),
    .B1(_04493_),
    .B2(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__mux2i_1 _10416_ (.A0(_04499_),
    .A1(_02983_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[23] ));
 sky130_fd_sc_hd__a21oi_1 _10417_ (.A1(\CPU_Xreg_value_a4[4][24] ),
    .A2(net29),
    .B1(net94),
    .Y(_04500_));
 sky130_fd_sc_hd__a22oi_1 _10418_ (.A1(\CPU_Xreg_value_a4[1][24] ),
    .A2(net36),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][24] ),
    .Y(_04501_));
 sky130_fd_sc_hd__a22oi_1 _10419_ (.A1(\CPU_Xreg_value_a4[8][24] ),
    .A2(net34),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][24] ),
    .Y(_04502_));
 sky130_fd_sc_hd__a22oi_1 _10420_ (.A1(\CPU_Xreg_value_a4[2][24] ),
    .A2(net33),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][24] ),
    .Y(_04503_));
 sky130_fd_sc_hd__nand4_2 _10421_ (.A(_04500_),
    .B(_04501_),
    .C(_04502_),
    .D(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__a22o_1 _10422_ (.A1(\CPU_Xreg_value_a4[3][24] ),
    .A2(net38),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][24] ),
    .X(_04505_));
 sky130_fd_sc_hd__a221oi_1 _10423_ (.A1(\CPU_Xreg_value_a4[6][24] ),
    .A2(_04258_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][24] ),
    .C1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__a22oi_1 _10424_ (.A1(\CPU_Xreg_value_a4[7][24] ),
    .A2(_04260_),
    .B1(net31),
    .B2(\CPU_Xreg_value_a4[12][24] ),
    .Y(_04507_));
 sky130_fd_sc_hd__a22oi_1 _10425_ (.A1(\CPU_Xreg_value_a4[15][24] ),
    .A2(_04268_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][24] ),
    .Y(_04508_));
 sky130_fd_sc_hd__nand3_1 _10426_ (.A(_04506_),
    .B(_04507_),
    .C(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__o22ai_4 _10427_ (.A1(net1542),
    .A2(_04231_),
    .B1(_04504_),
    .B2(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__and2_0 _10428_ (.A(_02997_),
    .B(_03007_),
    .X(_04511_));
 sky130_fd_sc_hd__mux2i_1 _10429_ (.A0(_04510_),
    .A1(_04511_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[24] ));
 sky130_fd_sc_hd__a21oi_1 _10430_ (.A1(\CPU_Xreg_value_a4[14][25] ),
    .A2(_04279_),
    .B1(net94),
    .Y(_04512_));
 sky130_fd_sc_hd__a22oi_1 _10431_ (.A1(\CPU_Xreg_value_a4[12][25] ),
    .A2(net31),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][25] ),
    .Y(_04513_));
 sky130_fd_sc_hd__a22oi_1 _10432_ (.A1(\CPU_Xreg_value_a4[6][25] ),
    .A2(_04258_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][25] ),
    .Y(_04514_));
 sky130_fd_sc_hd__a22oi_1 _10433_ (.A1(\CPU_Xreg_value_a4[10][25] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][25] ),
    .Y(_04515_));
 sky130_fd_sc_hd__nand4_1 _10434_ (.A(_04512_),
    .B(_04513_),
    .C(_04514_),
    .D(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__a22o_1 _10435_ (.A1(\CPU_Xreg_value_a4[2][25] ),
    .A2(net33),
    .B1(net29),
    .B2(\CPU_Xreg_value_a4[4][25] ),
    .X(_04517_));
 sky130_fd_sc_hd__a221oi_1 _10436_ (.A1(net1699),
    .A2(_04260_),
    .B1(net34),
    .B2(net1701),
    .C1(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a22oi_1 _10437_ (.A1(\CPU_Xreg_value_a4[11][25] ),
    .A2(_04275_),
    .B1(net40),
    .B2(net1703),
    .Y(_04519_));
 sky130_fd_sc_hd__a22oi_1 _10438_ (.A1(net1723),
    .A2(net36),
    .B1(_04281_),
    .B2(net1705),
    .Y(_04520_));
 sky130_fd_sc_hd__nand3_1 _10439_ (.A(_04518_),
    .B(_04519_),
    .C(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__o22ai_1 _10440_ (.A1(net1279),
    .A2(_04231_),
    .B1(_04516_),
    .B2(net1724),
    .Y(_04522_));
 sky130_fd_sc_hd__and2_0 _10441_ (.A(_03018_),
    .B(_03026_),
    .X(_04523_));
 sky130_fd_sc_hd__mux2i_1 _10442_ (.A0(net1725),
    .A1(_04523_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[25] ));
 sky130_fd_sc_hd__a21oi_1 _10443_ (.A1(\CPU_Xreg_value_a4[11][26] ),
    .A2(_04275_),
    .B1(net94),
    .Y(_04524_));
 sky130_fd_sc_hd__a22oi_1 _10444_ (.A1(\CPU_Xreg_value_a4[14][26] ),
    .A2(_04279_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][26] ),
    .Y(_04525_));
 sky130_fd_sc_hd__a22oi_1 _10445_ (.A1(\CPU_Xreg_value_a4[8][26] ),
    .A2(net34),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][26] ),
    .Y(_04526_));
 sky130_fd_sc_hd__a22oi_1 _10446_ (.A1(\CPU_Xreg_value_a4[1][26] ),
    .A2(net36),
    .B1(net31),
    .B2(\CPU_Xreg_value_a4[12][26] ),
    .Y(_04527_));
 sky130_fd_sc_hd__nand4_2 _10447_ (.A(_04524_),
    .B(_04525_),
    .C(_04526_),
    .D(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__a22o_1 _10448_ (.A1(\CPU_Xreg_value_a4[10][26] ),
    .A2(_04273_),
    .B1(net28),
    .B2(\CPU_Xreg_value_a4[4][26] ),
    .X(_04529_));
 sky130_fd_sc_hd__a221oi_1 _10449_ (.A1(\CPU_Xreg_value_a4[7][26] ),
    .A2(_04260_),
    .B1(net33),
    .B2(\CPU_Xreg_value_a4[2][26] ),
    .C1(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__a22oi_1 _10450_ (.A1(\CPU_Xreg_value_a4[6][26] ),
    .A2(_04258_),
    .B1(net38),
    .B2(\CPU_Xreg_value_a4[3][26] ),
    .Y(_04531_));
 sky130_fd_sc_hd__a22oi_1 _10451_ (.A1(\CPU_Xreg_value_a4[15][26] ),
    .A2(_04268_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][26] ),
    .Y(_04532_));
 sky130_fd_sc_hd__nand3_1 _10452_ (.A(_04530_),
    .B(_04531_),
    .C(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__o22ai_4 _10453_ (.A1(net1571),
    .A2(_04231_),
    .B1(_04528_),
    .B2(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3_1 _10454_ (.A(_03042_),
    .B(_03050_),
    .C(_03051_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_04535_),
    .B(_04292_),
    .Y(_04536_));
 sky130_fd_sc_hd__o21ai_0 _10456_ (.A1(_04292_),
    .A2(_04534_),
    .B1(_04536_),
    .Y(\CPU_src1_value_a2[26] ));
 sky130_fd_sc_hd__a21oi_1 _10457_ (.A1(\CPU_Xreg_value_a4[5][27] ),
    .A2(_04281_),
    .B1(net93),
    .Y(_04537_));
 sky130_fd_sc_hd__a22oi_1 _10458_ (.A1(\CPU_Xreg_value_a4[6][27] ),
    .A2(_04258_),
    .B1(_04260_),
    .B2(\CPU_Xreg_value_a4[7][27] ),
    .Y(_04538_));
 sky130_fd_sc_hd__a22oi_1 _10459_ (.A1(\CPU_Xreg_value_a4[10][27] ),
    .A2(_04273_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][27] ),
    .Y(_04539_));
 sky130_fd_sc_hd__a22oi_1 _10460_ (.A1(\CPU_Xreg_value_a4[12][27] ),
    .A2(net30),
    .B1(net27),
    .B2(\CPU_Xreg_value_a4[4][27] ),
    .Y(_04540_));
 sky130_fd_sc_hd__nand4_2 _10461_ (.A(_04537_),
    .B(_04538_),
    .C(_04539_),
    .D(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a22o_1 _10462_ (.A1(\CPU_Xreg_value_a4[2][27] ),
    .A2(net32),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][27] ),
    .X(_04542_));
 sky130_fd_sc_hd__a221oi_1 _10463_ (.A1(\CPU_Xreg_value_a4[11][27] ),
    .A2(_04275_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][27] ),
    .C1(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__a22oi_1 _10464_ (.A1(\CPU_Xreg_value_a4[8][27] ),
    .A2(net35),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][27] ),
    .Y(_04544_));
 sky130_fd_sc_hd__a22oi_1 _10465_ (.A1(\CPU_Xreg_value_a4[1][27] ),
    .A2(net36),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][27] ),
    .Y(_04545_));
 sky130_fd_sc_hd__nand3_1 _10466_ (.A(_04543_),
    .B(_04544_),
    .C(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__o22ai_4 _10467_ (.A1(net1848),
    .A2(_04231_),
    .B1(_04541_),
    .B2(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__mux2i_1 _10468_ (.A0(_04547_),
    .A1(_03074_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[27] ));
 sky130_fd_sc_hd__a21oi_1 _10469_ (.A1(\CPU_Xreg_value_a4[3][28] ),
    .A2(net38),
    .B1(net94),
    .Y(_04548_));
 sky130_fd_sc_hd__a22oi_1 _10470_ (.A1(\CPU_Xreg_value_a4[12][28] ),
    .A2(net30),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][28] ),
    .Y(_04549_));
 sky130_fd_sc_hd__a22oi_1 _10471_ (.A1(\CPU_Xreg_value_a4[15][28] ),
    .A2(_04268_),
    .B1(net28),
    .B2(\CPU_Xreg_value_a4[4][28] ),
    .Y(_04550_));
 sky130_fd_sc_hd__a22oi_1 _10472_ (.A1(\CPU_Xreg_value_a4[6][28] ),
    .A2(_04258_),
    .B1(net33),
    .B2(\CPU_Xreg_value_a4[2][28] ),
    .Y(_04551_));
 sky130_fd_sc_hd__nand4_1 _10473_ (.A(_04548_),
    .B(_04549_),
    .C(_04550_),
    .D(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a22o_1 _10474_ (.A1(\CPU_Xreg_value_a4[13][28] ),
    .A2(_04250_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][28] ),
    .X(_04553_));
 sky130_fd_sc_hd__a221oi_1 _10475_ (.A1(\CPU_Xreg_value_a4[1][28] ),
    .A2(net36),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][28] ),
    .C1(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__a22oi_1 _10476_ (.A1(\CPU_Xreg_value_a4[8][28] ),
    .A2(net34),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][28] ),
    .Y(_04555_));
 sky130_fd_sc_hd__a22oi_1 _10477_ (.A1(\CPU_Xreg_value_a4[7][28] ),
    .A2(_04260_),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][28] ),
    .Y(_04556_));
 sky130_fd_sc_hd__nand3_1 _10478_ (.A(_04554_),
    .B(_04555_),
    .C(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__o22ai_2 _10479_ (.A1(net1455),
    .A2(_04231_),
    .B1(_04552_),
    .B2(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__mux2i_1 _10480_ (.A0(_04558_),
    .A1(_03098_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[28] ));
 sky130_fd_sc_hd__a21o_1 _10481_ (.A1(net98),
    .A2(_03117_),
    .B1(_03135_),
    .X(_04559_));
 sky130_fd_sc_hd__a21oi_1 _10482_ (.A1(\CPU_Xreg_value_a4[4][29] ),
    .A2(net29),
    .B1(net94),
    .Y(_04560_));
 sky130_fd_sc_hd__a22oi_1 _10483_ (.A1(\CPU_Xreg_value_a4[2][29] ),
    .A2(net33),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][29] ),
    .Y(_04561_));
 sky130_fd_sc_hd__a22oi_1 _10484_ (.A1(\CPU_Xreg_value_a4[6][29] ),
    .A2(_04258_),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][29] ),
    .Y(_04562_));
 sky130_fd_sc_hd__a22oi_1 _10485_ (.A1(\CPU_Xreg_value_a4[15][29] ),
    .A2(_04268_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][29] ),
    .Y(_04563_));
 sky130_fd_sc_hd__nand4_1 _10486_ (.A(_04560_),
    .B(_04561_),
    .C(_04562_),
    .D(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__a22o_1 _10487_ (.A1(\CPU_Xreg_value_a4[1][29] ),
    .A2(net36),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][29] ),
    .X(_04565_));
 sky130_fd_sc_hd__a221oi_1 _10488_ (.A1(\CPU_Xreg_value_a4[12][29] ),
    .A2(net31),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][29] ),
    .C1(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__a22oi_1 _10489_ (.A1(\CPU_Xreg_value_a4[8][29] ),
    .A2(_04245_),
    .B1(net40),
    .B2(\CPU_Xreg_value_a4[3][29] ),
    .Y(_04567_));
 sky130_fd_sc_hd__a22oi_1 _10490_ (.A1(\CPU_Xreg_value_a4[7][29] ),
    .A2(_04260_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][29] ),
    .Y(_04568_));
 sky130_fd_sc_hd__nand3_1 _10491_ (.A(_04566_),
    .B(_04567_),
    .C(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__o22ai_1 _10492_ (.A1(net1266),
    .A2(_04231_),
    .B1(_04564_),
    .B2(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor2_1 _10493_ (.A(_04292_),
    .B(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21o_1 _10494_ (.A1(_04559_),
    .A2(_04292_),
    .B1(_04571_),
    .X(\CPU_src1_value_a2[29] ));
 sky130_fd_sc_hd__a21oi_1 _10495_ (.A1(\CPU_Xreg_value_a4[12][2] ),
    .A2(_04266_),
    .B1(net95),
    .Y(_04572_));
 sky130_fd_sc_hd__a22oi_1 _10496_ (.A1(\CPU_Xreg_value_a4[7][2] ),
    .A2(_04260_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][2] ),
    .Y(_04573_));
 sky130_fd_sc_hd__a22oi_1 _10497_ (.A1(\CPU_Xreg_value_a4[6][2] ),
    .A2(_04258_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][2] ),
    .Y(_04574_));
 sky130_fd_sc_hd__a22oi_1 _10498_ (.A1(\CPU_Xreg_value_a4[15][2] ),
    .A2(_04268_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][2] ),
    .Y(_04575_));
 sky130_fd_sc_hd__nand4_1 _10499_ (.A(_04572_),
    .B(_04573_),
    .C(_04574_),
    .D(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__a22o_1 _10500_ (.A1(\CPU_Xreg_value_a4[8][2] ),
    .A2(net35),
    .B1(net32),
    .B2(\CPU_Xreg_value_a4[2][2] ),
    .X(_04577_));
 sky130_fd_sc_hd__a221oi_1 _10501_ (.A1(\CPU_Xreg_value_a4[1][2] ),
    .A2(_04241_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][2] ),
    .C1(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__a22oi_1 _10502_ (.A1(\CPU_Xreg_value_a4[10][2] ),
    .A2(_04273_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][2] ),
    .Y(_04579_));
 sky130_fd_sc_hd__a22oi_1 _10503_ (.A1(\CPU_Xreg_value_a4[14][2] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][2] ),
    .Y(_04580_));
 sky130_fd_sc_hd__nand3_1 _10504_ (.A(_04578_),
    .B(_04579_),
    .C(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o22ai_4 _10505_ (.A1(net1666),
    .A2(_04231_),
    .B1(_04576_),
    .B2(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_1 _10506_ (.A(\CPU_result_a3[2] ),
    .B(_04292_),
    .Y(_04583_));
 sky130_fd_sc_hd__o21ai_0 _10507_ (.A1(_04292_),
    .A2(_04582_),
    .B1(_04583_),
    .Y(\CPU_src1_value_a2[2] ));
 sky130_fd_sc_hd__a21oi_1 _10508_ (.A1(\CPU_Xreg_value_a4[4][30] ),
    .A2(net28),
    .B1(net94),
    .Y(_04584_));
 sky130_fd_sc_hd__a22oi_1 _10509_ (.A1(\CPU_Xreg_value_a4[8][30] ),
    .A2(net34),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][30] ),
    .Y(_04585_));
 sky130_fd_sc_hd__a22oi_1 _10510_ (.A1(\CPU_Xreg_value_a4[1][30] ),
    .A2(net36),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][30] ),
    .Y(_04586_));
 sky130_fd_sc_hd__a22oi_1 _10511_ (.A1(\CPU_Xreg_value_a4[11][30] ),
    .A2(_04275_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][30] ),
    .Y(_04587_));
 sky130_fd_sc_hd__nand4_2 _10512_ (.A(_04584_),
    .B(_04585_),
    .C(_04586_),
    .D(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__a22o_1 _10513_ (.A1(\CPU_Xreg_value_a4[2][30] ),
    .A2(net33),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][30] ),
    .X(_04589_));
 sky130_fd_sc_hd__a221oi_1 _10514_ (.A1(\CPU_Xreg_value_a4[10][30] ),
    .A2(_04273_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][30] ),
    .C1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a22oi_1 _10515_ (.A1(\CPU_Xreg_value_a4[6][30] ),
    .A2(_04258_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][30] ),
    .Y(_04591_));
 sky130_fd_sc_hd__a22oi_1 _10516_ (.A1(\CPU_Xreg_value_a4[7][30] ),
    .A2(_04260_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][30] ),
    .Y(_04592_));
 sky130_fd_sc_hd__nand3_1 _10517_ (.A(_04590_),
    .B(_04591_),
    .C(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__o22ai_4 _10518_ (.A1(net1853),
    .A2(_04231_),
    .B1(_04588_),
    .B2(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__mux2i_1 _10519_ (.A0(_04594_),
    .A1(_03161_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[30] ));
 sky130_fd_sc_hd__a21oi_1 _10520_ (.A1(\CPU_Xreg_value_a4[15][31] ),
    .A2(_04268_),
    .B1(net93),
    .Y(_04595_));
 sky130_fd_sc_hd__a22oi_1 _10521_ (.A1(\CPU_Xreg_value_a4[14][31] ),
    .A2(_04279_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][31] ),
    .Y(_04596_));
 sky130_fd_sc_hd__a22oi_1 _10522_ (.A1(\CPU_Xreg_value_a4[10][31] ),
    .A2(_04273_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][31] ),
    .Y(_04597_));
 sky130_fd_sc_hd__a22oi_1 _10523_ (.A1(\CPU_Xreg_value_a4[6][31] ),
    .A2(_04258_),
    .B1(net32),
    .B2(\CPU_Xreg_value_a4[2][31] ),
    .Y(_04598_));
 sky130_fd_sc_hd__nand4_2 _10524_ (.A(_04595_),
    .B(_04596_),
    .C(_04597_),
    .D(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a22o_1 _10525_ (.A1(\CPU_Xreg_value_a4[1][31] ),
    .A2(net37),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][31] ),
    .X(_04600_));
 sky130_fd_sc_hd__a221oi_1 _10526_ (.A1(\CPU_Xreg_value_a4[4][31] ),
    .A2(net27),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][31] ),
    .C1(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__a22oi_1 _10527_ (.A1(\CPU_Xreg_value_a4[8][31] ),
    .A2(net34),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][31] ),
    .Y(_04602_));
 sky130_fd_sc_hd__a22oi_1 _10528_ (.A1(\CPU_Xreg_value_a4[7][31] ),
    .A2(_04260_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][31] ),
    .Y(_04603_));
 sky130_fd_sc_hd__nand3_1 _10529_ (.A(_04601_),
    .B(_04602_),
    .C(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__o22ai_4 _10530_ (.A1(net1683),
    .A2(_04231_),
    .B1(_04599_),
    .B2(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__mux2i_1 _10531_ (.A0(_04605_),
    .A1(_03189_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[31] ));
 sky130_fd_sc_hd__a21oi_1 _10532_ (.A1(\CPU_Xreg_value_a4[12][3] ),
    .A2(_04266_),
    .B1(net95),
    .Y(_04606_));
 sky130_fd_sc_hd__a22oi_1 _10533_ (.A1(\CPU_Xreg_value_a4[9][3] ),
    .A2(_04252_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][3] ),
    .Y(_04607_));
 sky130_fd_sc_hd__a22oi_1 _10534_ (.A1(\CPU_Xreg_value_a4[6][3] ),
    .A2(_04258_),
    .B1(net35),
    .B2(\CPU_Xreg_value_a4[8][3] ),
    .Y(_04608_));
 sky130_fd_sc_hd__a22oi_1 _10535_ (.A1(\CPU_Xreg_value_a4[15][3] ),
    .A2(_04268_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][3] ),
    .Y(_04609_));
 sky130_fd_sc_hd__nand4_1 _10536_ (.A(_04606_),
    .B(_04607_),
    .C(_04608_),
    .D(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__a22o_1 _10537_ (.A1(\CPU_Xreg_value_a4[1][3] ),
    .A2(_04241_),
    .B1(_04264_),
    .B2(\CPU_Xreg_value_a4[2][3] ),
    .X(_04611_));
 sky130_fd_sc_hd__a221oi_1 _10538_ (.A1(\CPU_Xreg_value_a4[7][3] ),
    .A2(_04260_),
    .B1(_04273_),
    .B2(\CPU_Xreg_value_a4[10][3] ),
    .C1(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__a22oi_1 _10539_ (.A1(\CPU_Xreg_value_a4[11][3] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][3] ),
    .Y(_04613_));
 sky130_fd_sc_hd__a22oi_1 _10540_ (.A1(\CPU_Xreg_value_a4[4][3] ),
    .A2(_04269_),
    .B1(_04234_),
    .B2(\CPU_Xreg_value_a4[3][3] ),
    .Y(_04614_));
 sky130_fd_sc_hd__nand3_1 _10541_ (.A(_04612_),
    .B(_04613_),
    .C(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__o22ai_4 _10542_ (.A1(net1520),
    .A2(_04231_),
    .B1(_04610_),
    .B2(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _10543_ (.A(\CPU_result_a3[3] ),
    .B(_04292_),
    .Y(_04617_));
 sky130_fd_sc_hd__o21ai_0 _10544_ (.A1(_04292_),
    .A2(_04616_),
    .B1(_04617_),
    .Y(\CPU_src1_value_a2[3] ));
 sky130_fd_sc_hd__a21oi_1 _10545_ (.A1(\CPU_Xreg_value_a4[3][4] ),
    .A2(net39),
    .B1(net95),
    .Y(_04618_));
 sky130_fd_sc_hd__a22oi_1 _10546_ (.A1(\CPU_Xreg_value_a4[9][4] ),
    .A2(_04252_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][4] ),
    .Y(_04619_));
 sky130_fd_sc_hd__a22oi_1 _10547_ (.A1(\CPU_Xreg_value_a4[6][4] ),
    .A2(_04258_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][4] ),
    .Y(_04620_));
 sky130_fd_sc_hd__a22oi_1 _10548_ (.A1(\CPU_Xreg_value_a4[11][4] ),
    .A2(_04275_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][4] ),
    .Y(_04621_));
 sky130_fd_sc_hd__nand4_2 _10549_ (.A(_04618_),
    .B(_04619_),
    .C(_04620_),
    .D(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__a22o_1 _10550_ (.A1(\CPU_Xreg_value_a4[12][4] ),
    .A2(net30),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][4] ),
    .X(_04623_));
 sky130_fd_sc_hd__a221oi_1 _10551_ (.A1(\CPU_Xreg_value_a4[7][4] ),
    .A2(_04260_),
    .B1(net35),
    .B2(\CPU_Xreg_value_a4[8][4] ),
    .C1(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__a22oi_1 _10552_ (.A1(\CPU_Xreg_value_a4[1][4] ),
    .A2(_04241_),
    .B1(net32),
    .B2(\CPU_Xreg_value_a4[2][4] ),
    .Y(_04625_));
 sky130_fd_sc_hd__a22oi_1 _10553_ (.A1(\CPU_Xreg_value_a4[10][4] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][4] ),
    .Y(_04626_));
 sky130_fd_sc_hd__nand3_1 _10554_ (.A(_04624_),
    .B(_04625_),
    .C(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__o22ai_4 _10555_ (.A1(net1849),
    .A2(_04231_),
    .B1(_04622_),
    .B2(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(\CPU_result_a3[4] ),
    .B(_04292_),
    .Y(_04629_));
 sky130_fd_sc_hd__o21ai_0 _10557_ (.A1(_04292_),
    .A2(_04628_),
    .B1(_04629_),
    .Y(\CPU_src1_value_a2[4] ));
 sky130_fd_sc_hd__a22oi_1 _10558_ (.A1(\CPU_Xreg_value_a4[6][5] ),
    .A2(_04258_),
    .B1(net32),
    .B2(\CPU_Xreg_value_a4[2][5] ),
    .Y(_04630_));
 sky130_fd_sc_hd__a22oi_1 _10559_ (.A1(\CPU_Xreg_value_a4[13][5] ),
    .A2(_04250_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][5] ),
    .Y(_04631_));
 sky130_fd_sc_hd__a22o_1 _10560_ (.A1(\CPU_Xreg_value_a4[15][5] ),
    .A2(_04268_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][5] ),
    .X(_04632_));
 sky130_fd_sc_hd__a221oi_1 _10561_ (.A1(\CPU_Xreg_value_a4[1][5] ),
    .A2(_04241_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][5] ),
    .C1(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__mux2i_1 _10562_ (.A0(\CPU_Xreg_value_a4[4][5] ),
    .A1(\CPU_Xreg_value_a4[12][5] ),
    .S(\CPU_rf_rd_index1_a2[3] ),
    .Y(_04634_));
 sky130_fd_sc_hd__o21ai_0 _10563_ (.A1(\CPU_Xreg_value_a4[8][5] ),
    .A2(_04244_),
    .B1(_04230_),
    .Y(_04635_));
 sky130_fd_sc_hd__a21oi_1 _10564_ (.A1(\CPU_rf_rd_index1_a2[2] ),
    .A2(_04634_),
    .B1(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__a221o_1 _10565_ (.A1(\CPU_Xreg_value_a4[10][5] ),
    .A2(_04273_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][5] ),
    .C1(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a221oi_1 _10566_ (.A1(\CPU_Xreg_value_a4[7][5] ),
    .A2(_04260_),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][5] ),
    .C1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand4_1 _10567_ (.A(_04630_),
    .B(_04631_),
    .C(_04633_),
    .D(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o21ai_2 _10568_ (.A1(net1618),
    .A2(_04231_),
    .B1(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__mux2i_1 _10569_ (.A0(_04640_),
    .A1(_03217_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[5] ));
 sky130_fd_sc_hd__a21oi_1 _10570_ (.A1(\CPU_Xreg_value_a4[4][6] ),
    .A2(net27),
    .B1(net93),
    .Y(_04641_));
 sky130_fd_sc_hd__a22oi_1 _10571_ (.A1(\CPU_Xreg_value_a4[10][6] ),
    .A2(_04273_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][6] ),
    .Y(_04642_));
 sky130_fd_sc_hd__a22oi_1 _10572_ (.A1(\CPU_Xreg_value_a4[6][6] ),
    .A2(_04258_),
    .B1(net30),
    .B2(\CPU_Xreg_value_a4[12][6] ),
    .Y(_04643_));
 sky130_fd_sc_hd__a22oi_1 _10573_ (.A1(\CPU_Xreg_value_a4[2][6] ),
    .A2(net32),
    .B1(_04279_),
    .B2(\CPU_Xreg_value_a4[14][6] ),
    .Y(_04644_));
 sky130_fd_sc_hd__nand4_2 _10574_ (.A(_04641_),
    .B(_04642_),
    .C(_04643_),
    .D(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__a22oi_1 _10575_ (.A1(\CPU_Xreg_value_a4[15][6] ),
    .A2(_04268_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][6] ),
    .Y(_04646_));
 sky130_fd_sc_hd__a22oi_1 _10576_ (.A1(\CPU_Xreg_value_a4[1][6] ),
    .A2(net36),
    .B1(_04260_),
    .B2(\CPU_Xreg_value_a4[7][6] ),
    .Y(_04647_));
 sky130_fd_sc_hd__a22o_1 _10577_ (.A1(\CPU_Xreg_value_a4[11][6] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][6] ),
    .X(_04648_));
 sky130_fd_sc_hd__a221oi_1 _10578_ (.A1(\CPU_Xreg_value_a4[8][6] ),
    .A2(net35),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][6] ),
    .C1(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand3_1 _10579_ (.A(_04646_),
    .B(_04647_),
    .C(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__o22ai_4 _10580_ (.A1(\CPU_Xreg_value_a4[0][6] ),
    .A2(_04231_),
    .B1(_04645_),
    .B2(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__mux2i_4 _10581_ (.A0(_04651_),
    .A1(_03225_),
    .S(_04292_),
    .Y(\CPU_src1_value_a2[6] ));
 sky130_fd_sc_hd__a21oi_1 _10582_ (.A1(\CPU_Xreg_value_a4[14][7] ),
    .A2(_04279_),
    .B1(net95),
    .Y(_04652_));
 sky130_fd_sc_hd__a22oi_1 _10583_ (.A1(\CPU_Xreg_value_a4[10][7] ),
    .A2(_04273_),
    .B1(_04264_),
    .B2(\CPU_Xreg_value_a4[2][7] ),
    .Y(_04653_));
 sky130_fd_sc_hd__a22oi_1 _10584_ (.A1(\CPU_Xreg_value_a4[1][7] ),
    .A2(_04241_),
    .B1(_04266_),
    .B2(\CPU_Xreg_value_a4[12][7] ),
    .Y(_04654_));
 sky130_fd_sc_hd__a22oi_1 _10585_ (.A1(\CPU_Xreg_value_a4[7][7] ),
    .A2(_04260_),
    .B1(net35),
    .B2(\CPU_Xreg_value_a4[8][7] ),
    .Y(_04655_));
 sky130_fd_sc_hd__nand4_1 _10586_ (.A(_04652_),
    .B(_04653_),
    .C(_04654_),
    .D(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__a22o_1 _10587_ (.A1(\CPU_Xreg_value_a4[6][7] ),
    .A2(_04258_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][7] ),
    .X(_04657_));
 sky130_fd_sc_hd__a221oi_1 _10588_ (.A1(\CPU_Xreg_value_a4[15][7] ),
    .A2(_04268_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][7] ),
    .C1(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__a22oi_1 _10589_ (.A1(\CPU_Xreg_value_a4[13][7] ),
    .A2(_04250_),
    .B1(_04234_),
    .B2(\CPU_Xreg_value_a4[3][7] ),
    .Y(_04659_));
 sky130_fd_sc_hd__a22oi_1 _10590_ (.A1(\CPU_Xreg_value_a4[11][7] ),
    .A2(_04275_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][7] ),
    .Y(_04660_));
 sky130_fd_sc_hd__nand3_1 _10591_ (.A(_04658_),
    .B(_04659_),
    .C(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__o22ai_4 _10592_ (.A1(\CPU_Xreg_value_a4[0][7] ),
    .A2(_04231_),
    .B1(_04656_),
    .B2(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand2_1 _10593_ (.A(_03235_),
    .B(_04292_),
    .Y(_04663_));
 sky130_fd_sc_hd__o21ai_0 _10594_ (.A1(_04292_),
    .A2(_04662_),
    .B1(_04663_),
    .Y(\CPU_src1_value_a2[7] ));
 sky130_fd_sc_hd__a21oi_1 _10595_ (.A1(\CPU_Xreg_value_a4[1][8] ),
    .A2(_04241_),
    .B1(net95),
    .Y(_04664_));
 sky130_fd_sc_hd__a22oi_1 _10596_ (.A1(\CPU_Xreg_value_a4[10][8] ),
    .A2(_04273_),
    .B1(_04268_),
    .B2(\CPU_Xreg_value_a4[15][8] ),
    .Y(_04665_));
 sky130_fd_sc_hd__a22oi_1 _10597_ (.A1(\CPU_Xreg_value_a4[11][8] ),
    .A2(_04275_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][8] ),
    .Y(_04666_));
 sky130_fd_sc_hd__a22oi_1 _10598_ (.A1(\CPU_Xreg_value_a4[14][8] ),
    .A2(_04279_),
    .B1(net39),
    .B2(\CPU_Xreg_value_a4[3][8] ),
    .Y(_04667_));
 sky130_fd_sc_hd__nand4_2 _10599_ (.A(_04664_),
    .B(_04665_),
    .C(_04666_),
    .D(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__a22o_1 _10600_ (.A1(\CPU_Xreg_value_a4[2][8] ),
    .A2(net32),
    .B1(_04266_),
    .B2(\CPU_Xreg_value_a4[12][8] ),
    .X(_04669_));
 sky130_fd_sc_hd__a221oi_1 _10601_ (.A1(\CPU_Xreg_value_a4[8][8] ),
    .A2(net35),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][8] ),
    .C1(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__a22oi_1 _10602_ (.A1(\CPU_Xreg_value_a4[6][8] ),
    .A2(_04258_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][8] ),
    .Y(_04671_));
 sky130_fd_sc_hd__a22oi_1 _10603_ (.A1(\CPU_Xreg_value_a4[7][8] ),
    .A2(_04260_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][8] ),
    .Y(_04672_));
 sky130_fd_sc_hd__nand3_1 _10604_ (.A(_04670_),
    .B(_04671_),
    .C(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__o22ai_4 _10605_ (.A1(net1850),
    .A2(_04231_),
    .B1(_04668_),
    .B2(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _10606_ (.A(_03248_),
    .B(_04292_),
    .Y(_04675_));
 sky130_fd_sc_hd__o21ai_0 _10607_ (.A1(_04292_),
    .A2(_04674_),
    .B1(_04675_),
    .Y(\CPU_src1_value_a2[8] ));
 sky130_fd_sc_hd__a21oi_1 _10608_ (.A1(\CPU_Xreg_value_a4[3][9] ),
    .A2(_04234_),
    .B1(net95),
    .Y(_04676_));
 sky130_fd_sc_hd__a22oi_1 _10609_ (.A1(\CPU_Xreg_value_a4[7][9] ),
    .A2(_04260_),
    .B1(_04266_),
    .B2(\CPU_Xreg_value_a4[12][9] ),
    .Y(_04677_));
 sky130_fd_sc_hd__a22oi_1 _10610_ (.A1(\CPU_Xreg_value_a4[10][9] ),
    .A2(_04273_),
    .B1(_04269_),
    .B2(\CPU_Xreg_value_a4[4][9] ),
    .Y(_04678_));
 sky130_fd_sc_hd__a22oi_1 _10611_ (.A1(\CPU_Xreg_value_a4[14][9] ),
    .A2(_04279_),
    .B1(_04252_),
    .B2(\CPU_Xreg_value_a4[9][9] ),
    .Y(_04679_));
 sky130_fd_sc_hd__nand4_1 _10612_ (.A(_04676_),
    .B(_04677_),
    .C(_04678_),
    .D(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__a22o_1 _10613_ (.A1(\CPU_Xreg_value_a4[1][9] ),
    .A2(_04241_),
    .B1(net35),
    .B2(\CPU_Xreg_value_a4[8][9] ),
    .X(_04681_));
 sky130_fd_sc_hd__a221oi_1 _10614_ (.A1(\CPU_Xreg_value_a4[2][9] ),
    .A2(_04264_),
    .B1(_04250_),
    .B2(\CPU_Xreg_value_a4[13][9] ),
    .C1(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__a22oi_1 _10615_ (.A1(\CPU_Xreg_value_a4[6][9] ),
    .A2(_04258_),
    .B1(_04275_),
    .B2(\CPU_Xreg_value_a4[11][9] ),
    .Y(_04683_));
 sky130_fd_sc_hd__a22oi_1 _10616_ (.A1(\CPU_Xreg_value_a4[15][9] ),
    .A2(_04268_),
    .B1(_04281_),
    .B2(\CPU_Xreg_value_a4[5][9] ),
    .Y(_04684_));
 sky130_fd_sc_hd__nand3_1 _10617_ (.A(_04682_),
    .B(_04683_),
    .C(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__o22ai_4 _10618_ (.A1(net1678),
    .A2(_04231_),
    .B1(_04680_),
    .B2(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _10619_ (.A(_03258_),
    .B(_04292_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21ai_0 _10620_ (.A1(_04292_),
    .A2(_04686_),
    .B1(_04687_),
    .Y(\CPU_src1_value_a2[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_102 ();
 sky130_fd_sc_hd__or4_4 _10625_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .C(\CPU_rf_rd_index2_a2[1] ),
    .D(\CPU_rf_rd_index2_a2[0] ),
    .X(_04692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_100 ();
 sky130_fd_sc_hd__nand2b_4 _10628_ (.A_N(\CPU_rf_rd_index2_a2[0] ),
    .B(\CPU_rf_rd_index2_a2[1] ),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_8 _10629_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .Y(_04696_));
 sky130_fd_sc_hd__nor2_8 _10630_ (.A(_04695_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_98 ();
 sky130_fd_sc_hd__nor4_4 _10633_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .C(\CPU_rf_rd_index2_a2[1] ),
    .D(\CPU_rf_rd_index2_a2[0] ),
    .Y(_04700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_97 ();
 sky130_fd_sc_hd__a21oi_1 _10635_ (.A1(\CPU_Xreg_value_a4[14][0] ),
    .A2(_04697_),
    .B1(net92),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2b_4 _10636_ (.A_N(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2_8 _10637_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .Y(_04704_));
 sky130_fd_sc_hd__nor2_8 _10638_ (.A(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_96 ();
 sky130_fd_sc_hd__nor3_4 _10640_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .C(_04696_),
    .Y(_04707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_95 ();
 sky130_fd_sc_hd__a22oi_1 _10642_ (.A1(\CPU_Xreg_value_a4[11][0] ),
    .A2(_04705_),
    .B1(net25),
    .B2(\CPU_Xreg_value_a4[12][0] ),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2b_4 _10643_ (.A_N(\CPU_rf_rd_index2_a2[1] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .Y(_04710_));
 sky130_fd_sc_hd__nor2_8 _10644_ (.A(_04703_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_94 ();
 sky130_fd_sc_hd__nor3_4 _10646_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .C(_04703_),
    .Y(_04713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_93 ();
 sky130_fd_sc_hd__a22oi_1 _10648_ (.A1(\CPU_Xreg_value_a4[9][0] ),
    .A2(_04711_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][0] ),
    .Y(_04715_));
 sky130_fd_sc_hd__nor3_4 _10649_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .C(_04695_),
    .Y(_04716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_92 ();
 sky130_fd_sc_hd__nand2b_4 _10651_ (.A_N(\CPU_rf_rd_index2_a2[3] ),
    .B(\CPU_rf_rd_index2_a2[2] ),
    .Y(_04718_));
 sky130_fd_sc_hd__nor2_8 _10652_ (.A(_04704_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__a22oi_1 _10655_ (.A1(\CPU_Xreg_value_a4[2][0] ),
    .A2(net20),
    .B1(_04719_),
    .B2(\CPU_Xreg_value_a4[7][0] ),
    .Y(_04722_));
 sky130_fd_sc_hd__nand4_2 _10656_ (.A(_04702_),
    .B(_04709_),
    .C(_04715_),
    .D(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nor3_4 _10657_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .C(_04704_),
    .Y(_04724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_89 ();
 sky130_fd_sc_hd__nor3_4 _10659_ (.A(\CPU_rf_rd_index2_a2[2] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .C(_04710_),
    .Y(_04726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_87 ();
 sky130_fd_sc_hd__nor2_8 _10662_ (.A(_04704_),
    .B(_04696_),
    .Y(_04729_));
 sky130_fd_sc_hd__nor2_8 _10663_ (.A(_04718_),
    .B(_04710_),
    .Y(_04730_));
 sky130_fd_sc_hd__a22o_1 _10664_ (.A1(\CPU_Xreg_value_a4[15][0] ),
    .A2(_04729_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][0] ),
    .X(_04731_));
 sky130_fd_sc_hd__a221oi_1 _10665_ (.A1(\CPU_Xreg_value_a4[3][0] ),
    .A2(net19),
    .B1(net17),
    .B2(\CPU_Xreg_value_a4[1][0] ),
    .C1(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__nor2_8 _10666_ (.A(_04703_),
    .B(_04695_),
    .Y(_04733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_85 ();
 sky130_fd_sc_hd__nor2_8 _10669_ (.A(_04696_),
    .B(_04710_),
    .Y(_04736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_83 ();
 sky130_fd_sc_hd__a22oi_1 _10672_ (.A1(\CPU_Xreg_value_a4[10][0] ),
    .A2(_04733_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][0] ),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_8 _10673_ (.A(_04695_),
    .B(_04718_),
    .Y(_04740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_82 ();
 sky130_fd_sc_hd__nor3_4 _10675_ (.A(\CPU_rf_rd_index2_a2[1] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .C(_04718_),
    .Y(_04742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_81 ();
 sky130_fd_sc_hd__a22oi_1 _10677_ (.A1(\CPU_Xreg_value_a4[6][0] ),
    .A2(_04740_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][0] ),
    .Y(_04744_));
 sky130_fd_sc_hd__nand3_1 _10678_ (.A(_04732_),
    .B(_04739_),
    .C(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__o22ai_4 _10679_ (.A1(\CPU_Xreg_value_a4[0][0] ),
    .A2(_04692_),
    .B1(_04723_),
    .B2(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__xnor2_1 _10680_ (.A(\CPU_rd_a3[0] ),
    .B(\CPU_rf_rd_index2_a2[0] ),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_1 _10681_ (.A(\CPU_rd_a3[3] ),
    .B(\CPU_rf_rd_index2_a2[3] ),
    .Y(_04748_));
 sky130_fd_sc_hd__xnor2_1 _10682_ (.A(\CPU_rd_a3[1] ),
    .B(\CPU_rf_rd_index2_a2[1] ),
    .Y(_04749_));
 sky130_fd_sc_hd__xnor2_1 _10683_ (.A(\CPU_rd_a3[2] ),
    .B(\CPU_rf_rd_index2_a2[2] ),
    .Y(_04750_));
 sky130_fd_sc_hd__nand4_2 _10684_ (.A(_04747_),
    .B(_04748_),
    .C(_04749_),
    .D(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nor2_8 _10685_ (.A(_04286_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_80 ();
 sky130_fd_sc_hd__mux2i_2 _10687_ (.A0(_04746_),
    .A1(_02560_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[0] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__a21oi_1 _10691_ (.A1(\CPU_Xreg_value_a4[7][10] ),
    .A2(_04719_),
    .B1(net91),
    .Y(_04757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__a22oi_1 _10694_ (.A1(\CPU_Xreg_value_a4[11][10] ),
    .A2(_04705_),
    .B1(net16),
    .B2(\CPU_Xreg_value_a4[1][10] ),
    .Y(_04760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_73 ();
 sky130_fd_sc_hd__a22oi_1 _10697_ (.A1(\CPU_Xreg_value_a4[5][10] ),
    .A2(_04730_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][10] ),
    .Y(_04763_));
 sky130_fd_sc_hd__a22oi_1 _10698_ (.A1(\CPU_Xreg_value_a4[10][10] ),
    .A2(_04733_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][10] ),
    .Y(_04764_));
 sky130_fd_sc_hd__nand4_1 _10699_ (.A(_04757_),
    .B(_04760_),
    .C(_04763_),
    .D(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_72 ();
 sky130_fd_sc_hd__a22o_1 _10701_ (.A1(\CPU_Xreg_value_a4[15][10] ),
    .A2(_04729_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][10] ),
    .X(_04767_));
 sky130_fd_sc_hd__a221oi_1 _10702_ (.A1(\CPU_Xreg_value_a4[2][10] ),
    .A2(net22),
    .B1(net18),
    .B2(\CPU_Xreg_value_a4[3][10] ),
    .C1(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__a22oi_1 _10703_ (.A1(\CPU_Xreg_value_a4[14][10] ),
    .A2(_04697_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][10] ),
    .Y(_04769_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_71 ();
 sky130_fd_sc_hd__a22oi_1 _10705_ (.A1(\CPU_Xreg_value_a4[12][10] ),
    .A2(net26),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][10] ),
    .Y(_04771_));
 sky130_fd_sc_hd__nand3_1 _10706_ (.A(_04768_),
    .B(_04769_),
    .C(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__o22ai_1 _10707_ (.A1(net1292),
    .A2(_04692_),
    .B1(_04765_),
    .B2(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__nand2_1 _10709_ (.A(_02635_),
    .B(_04752_),
    .Y(_04775_));
 sky130_fd_sc_hd__o21ai_0 _10710_ (.A1(_04752_),
    .A2(_04773_),
    .B1(_04775_),
    .Y(\CPU_src2_value_a2[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__a21oi_1 _10712_ (.A1(\CPU_Xreg_value_a4[9][11] ),
    .A2(_04711_),
    .B1(net90),
    .Y(_04777_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__a22oi_1 _10714_ (.A1(\CPU_Xreg_value_a4[5][11] ),
    .A2(_04730_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][11] ),
    .Y(_04779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_67 ();
 sky130_fd_sc_hd__a22oi_1 _10716_ (.A1(\CPU_Xreg_value_a4[11][11] ),
    .A2(_04705_),
    .B1(net19),
    .B2(\CPU_Xreg_value_a4[3][11] ),
    .Y(_04781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_66 ();
 sky130_fd_sc_hd__a22oi_1 _10718_ (.A1(\CPU_Xreg_value_a4[10][11] ),
    .A2(_04733_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][11] ),
    .Y(_04783_));
 sky130_fd_sc_hd__nand4_2 _10719_ (.A(_04777_),
    .B(_04779_),
    .C(_04781_),
    .D(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__a22o_1 _10722_ (.A1(\CPU_Xreg_value_a4[7][11] ),
    .A2(_04719_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][11] ),
    .X(_04787_));
 sky130_fd_sc_hd__a221oi_1 _10723_ (.A1(\CPU_Xreg_value_a4[2][11] ),
    .A2(net22),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][11] ),
    .C1(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__a22oi_1 _10724_ (.A1(\CPU_Xreg_value_a4[12][11] ),
    .A2(net26),
    .B1(net16),
    .B2(\CPU_Xreg_value_a4[1][11] ),
    .Y(_04789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__a22oi_1 _10727_ (.A1(\CPU_Xreg_value_a4[15][11] ),
    .A2(_04729_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][11] ),
    .Y(_04792_));
 sky130_fd_sc_hd__nand3_1 _10728_ (.A(_04788_),
    .B(_04789_),
    .C(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__o22ai_4 _10729_ (.A1(net1504),
    .A2(_04692_),
    .B1(_04784_),
    .B2(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _10730_ (.A(_04338_),
    .B(_04752_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ai_0 _10731_ (.A1(_04752_),
    .A2(_04794_),
    .B1(_04795_),
    .Y(\CPU_src2_value_a2[11] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__a21oi_1 _10734_ (.A1(\CPU_Xreg_value_a4[1][12] ),
    .A2(_04726_),
    .B1(_04700_),
    .Y(_04798_));
 sky130_fd_sc_hd__a22oi_1 _10735_ (.A1(\CPU_Xreg_value_a4[10][12] ),
    .A2(_04733_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][12] ),
    .Y(_04799_));
 sky130_fd_sc_hd__a22oi_1 _10736_ (.A1(\CPU_Xreg_value_a4[9][12] ),
    .A2(_04711_),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][12] ),
    .Y(_04800_));
 sky130_fd_sc_hd__a22oi_1 _10737_ (.A1(\CPU_Xreg_value_a4[11][12] ),
    .A2(_04705_),
    .B1(_04724_),
    .B2(\CPU_Xreg_value_a4[3][12] ),
    .Y(_04801_));
 sky130_fd_sc_hd__nand4_1 _10738_ (.A(_04798_),
    .B(_04799_),
    .C(_04800_),
    .D(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__a22o_1 _10739_ (.A1(\CPU_Xreg_value_a4[2][12] ),
    .A2(_04716_),
    .B1(_04719_),
    .B2(\CPU_Xreg_value_a4[7][12] ),
    .X(_04803_));
 sky130_fd_sc_hd__a221oi_1 _10740_ (.A1(\CPU_Xreg_value_a4[12][12] ),
    .A2(_04707_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][12] ),
    .C1(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_58 ();
 sky130_fd_sc_hd__a22oi_1 _10743_ (.A1(\CPU_Xreg_value_a4[13][12] ),
    .A2(_04736_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][12] ),
    .Y(_04807_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_57 ();
 sky130_fd_sc_hd__a22oi_1 _10745_ (.A1(\CPU_Xreg_value_a4[15][12] ),
    .A2(_04729_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][12] ),
    .Y(_04809_));
 sky130_fd_sc_hd__nand3_1 _10746_ (.A(_04804_),
    .B(_04807_),
    .C(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__o22ai_4 _10747_ (.A1(\CPU_Xreg_value_a4[0][12] ),
    .A2(_04692_),
    .B1(_04802_),
    .B2(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(_02710_),
    .B(_04752_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21ai_0 _10749_ (.A1(_04752_),
    .A2(_04811_),
    .B1(_04812_),
    .Y(\CPU_src2_value_a2[12] ));
 sky130_fd_sc_hd__a21oi_1 _10750_ (.A1(\CPU_Xreg_value_a4[6][13] ),
    .A2(_04740_),
    .B1(net91),
    .Y(_04813_));
 sky130_fd_sc_hd__a22oi_1 _10751_ (.A1(\CPU_Xreg_value_a4[7][13] ),
    .A2(_04719_),
    .B1(net26),
    .B2(\CPU_Xreg_value_a4[12][13] ),
    .Y(_04814_));
 sky130_fd_sc_hd__a22oi_1 _10752_ (.A1(\CPU_Xreg_value_a4[13][13] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][13] ),
    .Y(_04815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_56 ();
 sky130_fd_sc_hd__a22oi_1 _10754_ (.A1(\CPU_Xreg_value_a4[10][13] ),
    .A2(_04733_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][13] ),
    .Y(_04817_));
 sky130_fd_sc_hd__nand4_1 _10755_ (.A(_04813_),
    .B(_04814_),
    .C(_04815_),
    .D(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__a22o_1 _10758_ (.A1(\CPU_Xreg_value_a4[15][13] ),
    .A2(_04729_),
    .B1(net16),
    .B2(\CPU_Xreg_value_a4[1][13] ),
    .X(_04821_));
 sky130_fd_sc_hd__a221oi_1 _10759_ (.A1(\CPU_Xreg_value_a4[11][13] ),
    .A2(_04705_),
    .B1(net18),
    .B2(\CPU_Xreg_value_a4[3][13] ),
    .C1(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__a22oi_1 _10760_ (.A1(\CPU_Xreg_value_a4[9][13] ),
    .A2(_04711_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][13] ),
    .Y(_04823_));
 sky130_fd_sc_hd__a22oi_1 _10761_ (.A1(\CPU_Xreg_value_a4[2][13] ),
    .A2(net22),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][13] ),
    .Y(_04824_));
 sky130_fd_sc_hd__nand3_1 _10762_ (.A(_04822_),
    .B(_04823_),
    .C(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__o22ai_4 _10763_ (.A1(net1503),
    .A2(_04692_),
    .B1(_04818_),
    .B2(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__mux2i_1 _10764_ (.A0(_04826_),
    .A1(_04369_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[13] ));
 sky130_fd_sc_hd__a21oi_1 _10765_ (.A1(\CPU_Xreg_value_a4[7][14] ),
    .A2(_04719_),
    .B1(net91),
    .Y(_04827_));
 sky130_fd_sc_hd__a22oi_1 _10766_ (.A1(\CPU_Xreg_value_a4[6][14] ),
    .A2(_04740_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][14] ),
    .Y(_04828_));
 sky130_fd_sc_hd__a22oi_1 _10767_ (.A1(\CPU_Xreg_value_a4[3][14] ),
    .A2(net18),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][14] ),
    .Y(_04829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__a22oi_1 _10769_ (.A1(\CPU_Xreg_value_a4[10][14] ),
    .A2(_04733_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][14] ),
    .Y(_04831_));
 sky130_fd_sc_hd__nand4_1 _10770_ (.A(_04827_),
    .B(_04828_),
    .C(_04829_),
    .D(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a22o_1 _10771_ (.A1(\CPU_Xreg_value_a4[1][14] ),
    .A2(net17),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][14] ),
    .X(_04833_));
 sky130_fd_sc_hd__a221oi_1 _10772_ (.A1(\CPU_Xreg_value_a4[2][14] ),
    .A2(net22),
    .B1(net26),
    .B2(net1744),
    .C1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__a22oi_1 _10773_ (.A1(\CPU_Xreg_value_a4[14][14] ),
    .A2(_04697_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][14] ),
    .Y(_04835_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__a22oi_1 _10775_ (.A1(\CPU_Xreg_value_a4[11][14] ),
    .A2(_04705_),
    .B1(_04711_),
    .B2(net1760),
    .Y(_04837_));
 sky130_fd_sc_hd__nand3_1 _10776_ (.A(_04834_),
    .B(_04835_),
    .C(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__o22ai_1 _10777_ (.A1(net1269),
    .A2(_04692_),
    .B1(_04832_),
    .B2(net1761),
    .Y(_04839_));
 sky130_fd_sc_hd__mux2i_1 _10778_ (.A0(net1762),
    .A1(_02764_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[14] ));
 sky130_fd_sc_hd__a21oi_1 _10779_ (.A1(\CPU_Xreg_value_a4[5][15] ),
    .A2(_04730_),
    .B1(_04700_),
    .Y(_04840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__a22oi_1 _10781_ (.A1(\CPU_Xreg_value_a4[12][15] ),
    .A2(net26),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][15] ),
    .Y(_04842_));
 sky130_fd_sc_hd__a22oi_1 _10782_ (.A1(\CPU_Xreg_value_a4[11][15] ),
    .A2(_04705_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][15] ),
    .Y(_04843_));
 sky130_fd_sc_hd__a22oi_1 _10783_ (.A1(\CPU_Xreg_value_a4[13][15] ),
    .A2(_04736_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][15] ),
    .Y(_04844_));
 sky130_fd_sc_hd__nand4_1 _10784_ (.A(_04840_),
    .B(_04842_),
    .C(_04843_),
    .D(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__a22o_1 _10785_ (.A1(\CPU_Xreg_value_a4[7][15] ),
    .A2(_04719_),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][15] ),
    .X(_04846_));
 sky130_fd_sc_hd__a221oi_1 _10786_ (.A1(\CPU_Xreg_value_a4[1][15] ),
    .A2(net17),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][15] ),
    .C1(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__a22oi_2 _10787_ (.A1(\CPU_Xreg_value_a4[2][15] ),
    .A2(net21),
    .B1(net19),
    .B2(\CPU_Xreg_value_a4[3][15] ),
    .Y(_04848_));
 sky130_fd_sc_hd__a22oi_1 _10788_ (.A1(\CPU_Xreg_value_a4[15][15] ),
    .A2(_04729_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][15] ),
    .Y(_04849_));
 sky130_fd_sc_hd__nand3_1 _10789_ (.A(_04847_),
    .B(_04848_),
    .C(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__o22ai_1 _10790_ (.A1(net1307),
    .A2(_04692_),
    .B1(_04845_),
    .B2(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(_02782_),
    .B(_04752_),
    .Y(_04852_));
 sky130_fd_sc_hd__o21ai_0 _10792_ (.A1(_04752_),
    .A2(_04851_),
    .B1(_04852_),
    .Y(\CPU_src2_value_a2[15] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__a21oi_1 _10794_ (.A1(net1424),
    .A2(_04730_),
    .B1(_04700_),
    .Y(_04854_));
 sky130_fd_sc_hd__a22oi_1 _10795_ (.A1(\CPU_Xreg_value_a4[7][16] ),
    .A2(_04719_),
    .B1(net18),
    .B2(net1384),
    .Y(_04855_));
 sky130_fd_sc_hd__a22oi_1 _10796_ (.A1(\CPU_Xreg_value_a4[15][16] ),
    .A2(_04729_),
    .B1(_04736_),
    .B2(net1737),
    .Y(_04856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__a22oi_1 _10798_ (.A1(\CPU_Xreg_value_a4[12][16] ),
    .A2(net26),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][16] ),
    .Y(_04858_));
 sky130_fd_sc_hd__nand4_1 _10799_ (.A(_04854_),
    .B(_04855_),
    .C(_04856_),
    .D(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__a22o_1 _10801_ (.A1(\CPU_Xreg_value_a4[6][16] ),
    .A2(_04740_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][16] ),
    .X(_04861_));
 sky130_fd_sc_hd__a221oi_1 _10802_ (.A1(net1439),
    .A2(net22),
    .B1(net17),
    .B2(net1442),
    .C1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__a22oi_1 _10803_ (.A1(\CPU_Xreg_value_a4[10][16] ),
    .A2(_04733_),
    .B1(_04711_),
    .B2(net1390),
    .Y(_04863_));
 sky130_fd_sc_hd__a22oi_1 _10804_ (.A1(\CPU_Xreg_value_a4[11][16] ),
    .A2(_04705_),
    .B1(_04713_),
    .B2(net1452),
    .Y(_04864_));
 sky130_fd_sc_hd__nand3_1 _10805_ (.A(_04862_),
    .B(_04863_),
    .C(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__o22ai_1 _10806_ (.A1(net1312),
    .A2(_04692_),
    .B1(_04859_),
    .B2(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__mux2i_1 _10807_ (.A0(_04866_),
    .A1(_02807_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[16] ));
 sky130_fd_sc_hd__a21oi_1 _10808_ (.A1(net1498),
    .A2(_04729_),
    .B1(_04700_),
    .Y(_04867_));
 sky130_fd_sc_hd__a22oi_1 _10809_ (.A1(\CPU_Xreg_value_a4[9][17] ),
    .A2(_04711_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][17] ),
    .Y(_04868_));
 sky130_fd_sc_hd__a22oi_1 _10810_ (.A1(\CPU_Xreg_value_a4[11][17] ),
    .A2(_04705_),
    .B1(net25),
    .B2(\CPU_Xreg_value_a4[12][17] ),
    .Y(_04869_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__a22oi_1 _10812_ (.A1(\CPU_Xreg_value_a4[7][17] ),
    .A2(_04719_),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][17] ),
    .Y(_04871_));
 sky130_fd_sc_hd__nand4_1 _10813_ (.A(_04867_),
    .B(_04868_),
    .C(_04869_),
    .D(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__a22o_1 _10814_ (.A1(\CPU_Xreg_value_a4[13][17] ),
    .A2(_04736_),
    .B1(net17),
    .B2(\CPU_Xreg_value_a4[1][17] ),
    .X(_04873_));
 sky130_fd_sc_hd__a221oi_1 _10815_ (.A1(\CPU_Xreg_value_a4[2][17] ),
    .A2(net20),
    .B1(net19),
    .B2(\CPU_Xreg_value_a4[3][17] ),
    .C1(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__a22oi_1 _10816_ (.A1(\CPU_Xreg_value_a4[6][17] ),
    .A2(_04740_),
    .B1(net15),
    .B2(net1526),
    .Y(_04875_));
 sky130_fd_sc_hd__a22oi_1 _10817_ (.A1(\CPU_Xreg_value_a4[5][17] ),
    .A2(_04730_),
    .B1(_04697_),
    .B2(net1794),
    .Y(_04876_));
 sky130_fd_sc_hd__nand3_1 _10818_ (.A(_04874_),
    .B(_04875_),
    .C(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__o22ai_2 _10819_ (.A1(net1418),
    .A2(_04692_),
    .B1(_04872_),
    .B2(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__mux2i_1 _10821_ (.A0(_04878_),
    .A1(_02832_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[17] ));
 sky130_fd_sc_hd__a21oi_1 _10822_ (.A1(\CPU_Xreg_value_a4[4][18] ),
    .A2(net15),
    .B1(net91),
    .Y(_04880_));
 sky130_fd_sc_hd__a22oi_1 _10823_ (.A1(\CPU_Xreg_value_a4[2][18] ),
    .A2(net22),
    .B1(_04719_),
    .B2(\CPU_Xreg_value_a4[7][18] ),
    .Y(_04881_));
 sky130_fd_sc_hd__a22oi_1 _10824_ (.A1(\CPU_Xreg_value_a4[11][18] ),
    .A2(_04705_),
    .B1(net26),
    .B2(\CPU_Xreg_value_a4[12][18] ),
    .Y(_04882_));
 sky130_fd_sc_hd__a22oi_1 _10825_ (.A1(\CPU_Xreg_value_a4[10][18] ),
    .A2(_04733_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][18] ),
    .Y(_04883_));
 sky130_fd_sc_hd__nand4_1 _10826_ (.A(_04880_),
    .B(_04881_),
    .C(_04882_),
    .D(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__a22oi_1 _10827_ (.A1(\CPU_Xreg_value_a4[1][18] ),
    .A2(net16),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][18] ),
    .Y(_04885_));
 sky130_fd_sc_hd__a22oi_1 _10828_ (.A1(\CPU_Xreg_value_a4[5][18] ),
    .A2(_04730_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][18] ),
    .Y(_04886_));
 sky130_fd_sc_hd__a22oi_1 _10829_ (.A1(\CPU_Xreg_value_a4[15][18] ),
    .A2(_04729_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][18] ),
    .Y(_04887_));
 sky130_fd_sc_hd__a22oi_1 _10830_ (.A1(\CPU_Xreg_value_a4[3][18] ),
    .A2(net18),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][18] ),
    .Y(_04888_));
 sky130_fd_sc_hd__nand4_1 _10831_ (.A(_04885_),
    .B(_04886_),
    .C(_04887_),
    .D(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__o22ai_2 _10832_ (.A1(net1610),
    .A2(_04692_),
    .B1(_04884_),
    .B2(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__mux2i_1 _10833_ (.A0(_04890_),
    .A1(_02853_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[18] ));
 sky130_fd_sc_hd__a21oi_1 _10834_ (.A1(\CPU_Xreg_value_a4[15][19] ),
    .A2(_04729_),
    .B1(_04700_),
    .Y(_04891_));
 sky130_fd_sc_hd__a22oi_1 _10835_ (.A1(\CPU_Xreg_value_a4[7][19] ),
    .A2(_04719_),
    .B1(net26),
    .B2(\CPU_Xreg_value_a4[12][19] ),
    .Y(_04892_));
 sky130_fd_sc_hd__a22oi_1 _10836_ (.A1(\CPU_Xreg_value_a4[8][19] ),
    .A2(net23),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][19] ),
    .Y(_04893_));
 sky130_fd_sc_hd__a22oi_1 _10837_ (.A1(\CPU_Xreg_value_a4[3][19] ),
    .A2(net18),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][19] ),
    .Y(_04894_));
 sky130_fd_sc_hd__nand4_1 _10838_ (.A(_04891_),
    .B(_04892_),
    .C(_04893_),
    .D(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__a22o_1 _10839_ (.A1(\CPU_Xreg_value_a4[1][19] ),
    .A2(net17),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][19] ),
    .X(_04896_));
 sky130_fd_sc_hd__a221oi_1 _10840_ (.A1(\CPU_Xreg_value_a4[11][19] ),
    .A2(_04705_),
    .B1(net20),
    .B2(\CPU_Xreg_value_a4[2][19] ),
    .C1(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__a22oi_1 _10841_ (.A1(\CPU_Xreg_value_a4[10][19] ),
    .A2(_04733_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][19] ),
    .Y(_04898_));
 sky130_fd_sc_hd__a22oi_1 _10842_ (.A1(\CPU_Xreg_value_a4[13][19] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][19] ),
    .Y(_04899_));
 sky130_fd_sc_hd__nand3_1 _10843_ (.A(_04897_),
    .B(_04898_),
    .C(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__o22ai_2 _10844_ (.A1(net1409),
    .A2(_04692_),
    .B1(_04895_),
    .B2(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21ai_0 _10845_ (.A1(_02866_),
    .A2(_02881_),
    .B1(_04752_),
    .Y(_04902_));
 sky130_fd_sc_hd__o21ai_0 _10846_ (.A1(_04752_),
    .A2(_04901_),
    .B1(_04902_),
    .Y(\CPU_src2_value_a2[19] ));
 sky130_fd_sc_hd__a21oi_1 _10847_ (.A1(\CPU_Xreg_value_a4[6][1] ),
    .A2(_04740_),
    .B1(net92),
    .Y(_04903_));
 sky130_fd_sc_hd__a22oi_1 _10848_ (.A1(\CPU_Xreg_value_a4[2][1] ),
    .A2(_04716_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][1] ),
    .Y(_04904_));
 sky130_fd_sc_hd__a22oi_1 _10849_ (.A1(\CPU_Xreg_value_a4[11][1] ),
    .A2(_04705_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][1] ),
    .Y(_04905_));
 sky130_fd_sc_hd__a22oi_1 _10850_ (.A1(\CPU_Xreg_value_a4[14][1] ),
    .A2(_04697_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][1] ),
    .Y(_04906_));
 sky130_fd_sc_hd__nand4_1 _10851_ (.A(_04903_),
    .B(_04904_),
    .C(_04905_),
    .D(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__a22o_1 _10852_ (.A1(\CPU_Xreg_value_a4[7][1] ),
    .A2(_04719_),
    .B1(_04726_),
    .B2(\CPU_Xreg_value_a4[1][1] ),
    .X(_04908_));
 sky130_fd_sc_hd__a221oi_1 _10853_ (.A1(\CPU_Xreg_value_a4[10][1] ),
    .A2(_04733_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][1] ),
    .C1(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a22oi_1 _10854_ (.A1(\CPU_Xreg_value_a4[3][1] ),
    .A2(_04724_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][1] ),
    .Y(_04910_));
 sky130_fd_sc_hd__a22oi_1 _10855_ (.A1(\CPU_Xreg_value_a4[12][1] ),
    .A2(_04707_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][1] ),
    .Y(_04911_));
 sky130_fd_sc_hd__nand3_1 _10856_ (.A(_04909_),
    .B(_04910_),
    .C(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__o22ai_4 _10857_ (.A1(net1854),
    .A2(_04692_),
    .B1(_04907_),
    .B2(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_1 _10858_ (.A(_02888_),
    .B(_04752_),
    .Y(_04914_));
 sky130_fd_sc_hd__o21ai_0 _10859_ (.A1(_04752_),
    .A2(_04913_),
    .B1(_04914_),
    .Y(\CPU_src2_value_a2[1] ));
 sky130_fd_sc_hd__a21oi_1 _10860_ (.A1(\CPU_Xreg_value_a4[5][20] ),
    .A2(_04730_),
    .B1(net92),
    .Y(_04915_));
 sky130_fd_sc_hd__a22oi_1 _10861_ (.A1(\CPU_Xreg_value_a4[12][20] ),
    .A2(net25),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][20] ),
    .Y(_04916_));
 sky130_fd_sc_hd__a22oi_1 _10862_ (.A1(\CPU_Xreg_value_a4[11][20] ),
    .A2(_04705_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][20] ),
    .Y(_04917_));
 sky130_fd_sc_hd__a22oi_1 _10863_ (.A1(\CPU_Xreg_value_a4[2][20] ),
    .A2(net20),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][20] ),
    .Y(_04918_));
 sky130_fd_sc_hd__nand4_1 _10864_ (.A(_04915_),
    .B(_04916_),
    .C(_04917_),
    .D(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a22o_1 _10865_ (.A1(\CPU_Xreg_value_a4[1][20] ),
    .A2(net17),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][20] ),
    .X(_04920_));
 sky130_fd_sc_hd__a221oi_1 _10866_ (.A1(\CPU_Xreg_value_a4[7][20] ),
    .A2(_04719_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][20] ),
    .C1(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__a22oi_1 _10867_ (.A1(\CPU_Xreg_value_a4[3][20] ),
    .A2(net19),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][20] ),
    .Y(_04922_));
 sky130_fd_sc_hd__a22oi_1 _10868_ (.A1(\CPU_Xreg_value_a4[10][20] ),
    .A2(_04733_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][20] ),
    .Y(_04923_));
 sky130_fd_sc_hd__nand3_1 _10869_ (.A(_04921_),
    .B(_04922_),
    .C(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__o22ai_4 _10870_ (.A1(net1675),
    .A2(_04692_),
    .B1(_04919_),
    .B2(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__mux2i_1 _10871_ (.A0(_04925_),
    .A1(_02908_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[20] ));
 sky130_fd_sc_hd__a21oi_1 _10872_ (.A1(\CPU_Xreg_value_a4[4][21] ),
    .A2(net14),
    .B1(net90),
    .Y(_04926_));
 sky130_fd_sc_hd__a22oi_1 _10873_ (.A1(\CPU_Xreg_value_a4[13][21] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][21] ),
    .Y(_04927_));
 sky130_fd_sc_hd__a22oi_1 _10874_ (.A1(\CPU_Xreg_value_a4[3][21] ),
    .A2(_04724_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][21] ),
    .Y(_04928_));
 sky130_fd_sc_hd__a22oi_1 _10875_ (.A1(\CPU_Xreg_value_a4[12][21] ),
    .A2(_04707_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][21] ),
    .Y(_04929_));
 sky130_fd_sc_hd__nand4_2 _10876_ (.A(_04926_),
    .B(_04927_),
    .C(_04928_),
    .D(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__a22o_1 _10877_ (.A1(\CPU_Xreg_value_a4[7][21] ),
    .A2(_04719_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][21] ),
    .X(_04931_));
 sky130_fd_sc_hd__a221oi_1 _10878_ (.A1(\CPU_Xreg_value_a4[2][21] ),
    .A2(net21),
    .B1(net17),
    .B2(\CPU_Xreg_value_a4[1][21] ),
    .C1(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__a22oi_1 _10879_ (.A1(\CPU_Xreg_value_a4[6][21] ),
    .A2(_04740_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][21] ),
    .Y(_04933_));
 sky130_fd_sc_hd__a22oi_1 _10880_ (.A1(\CPU_Xreg_value_a4[11][21] ),
    .A2(_04705_),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][21] ),
    .Y(_04934_));
 sky130_fd_sc_hd__nand3_1 _10881_ (.A(_04932_),
    .B(_04933_),
    .C(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__o22ai_4 _10882_ (.A1(net1671),
    .A2(_04692_),
    .B1(_04930_),
    .B2(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__mux2i_1 _10883_ (.A0(_04936_),
    .A1(_02934_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[21] ));
 sky130_fd_sc_hd__a21oi_1 _10884_ (.A1(\CPU_Xreg_value_a4[5][22] ),
    .A2(_04730_),
    .B1(net91),
    .Y(_04937_));
 sky130_fd_sc_hd__a22oi_1 _10885_ (.A1(\CPU_Xreg_value_a4[7][22] ),
    .A2(_04719_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][22] ),
    .Y(_04938_));
 sky130_fd_sc_hd__a22oi_1 _10886_ (.A1(\CPU_Xreg_value_a4[12][22] ),
    .A2(net26),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][22] ),
    .Y(_04939_));
 sky130_fd_sc_hd__a22oi_1 _10887_ (.A1(\CPU_Xreg_value_a4[10][22] ),
    .A2(_04733_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][22] ),
    .Y(_04940_));
 sky130_fd_sc_hd__nand4_1 _10888_ (.A(_04937_),
    .B(_04938_),
    .C(_04939_),
    .D(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__a22o_1 _10889_ (.A1(\CPU_Xreg_value_a4[1][22] ),
    .A2(net16),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][22] ),
    .X(_04942_));
 sky130_fd_sc_hd__a221oi_1 _10890_ (.A1(\CPU_Xreg_value_a4[2][22] ),
    .A2(net20),
    .B1(net18),
    .B2(\CPU_Xreg_value_a4[3][22] ),
    .C1(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__a22oi_1 _10891_ (.A1(\CPU_Xreg_value_a4[11][22] ),
    .A2(_04705_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][22] ),
    .Y(_04944_));
 sky130_fd_sc_hd__a22oi_1 _10892_ (.A1(\CPU_Xreg_value_a4[6][22] ),
    .A2(_04740_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][22] ),
    .Y(_04945_));
 sky130_fd_sc_hd__nand3_1 _10893_ (.A(_04943_),
    .B(_04944_),
    .C(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__o22ai_4 _10894_ (.A1(net1607),
    .A2(_04692_),
    .B1(_04941_),
    .B2(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__mux2i_1 _10895_ (.A0(_04947_),
    .A1(_02959_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[22] ));
 sky130_fd_sc_hd__a21oi_1 _10896_ (.A1(\CPU_Xreg_value_a4[4][23] ),
    .A2(net14),
    .B1(net90),
    .Y(_04948_));
 sky130_fd_sc_hd__a22oi_1 _10897_ (.A1(\CPU_Xreg_value_a4[3][23] ),
    .A2(net19),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][23] ),
    .Y(_04949_));
 sky130_fd_sc_hd__a22oi_1 _10898_ (.A1(\CPU_Xreg_value_a4[11][23] ),
    .A2(_04705_),
    .B1(net25),
    .B2(\CPU_Xreg_value_a4[12][23] ),
    .Y(_04950_));
 sky130_fd_sc_hd__a22oi_1 _10899_ (.A1(\CPU_Xreg_value_a4[15][23] ),
    .A2(_04729_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][23] ),
    .Y(_04951_));
 sky130_fd_sc_hd__nand4_1 _10900_ (.A(_04948_),
    .B(_04949_),
    .C(_04950_),
    .D(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__a22o_1 _10901_ (.A1(\CPU_Xreg_value_a4[9][23] ),
    .A2(_04711_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][23] ),
    .X(_04953_));
 sky130_fd_sc_hd__a221oi_1 _10902_ (.A1(\CPU_Xreg_value_a4[2][23] ),
    .A2(net21),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][23] ),
    .C1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a22oi_1 _10903_ (.A1(\CPU_Xreg_value_a4[1][23] ),
    .A2(net17),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][23] ),
    .Y(_04955_));
 sky130_fd_sc_hd__a22oi_1 _10904_ (.A1(\CPU_Xreg_value_a4[7][23] ),
    .A2(_04719_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][23] ),
    .Y(_04956_));
 sky130_fd_sc_hd__nand3_1 _10905_ (.A(_04954_),
    .B(_04955_),
    .C(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__o22ai_4 _10906_ (.A1(net1511),
    .A2(_04692_),
    .B1(_04952_),
    .B2(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__mux2i_1 _10907_ (.A0(_04958_),
    .A1(_02983_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[23] ));
 sky130_fd_sc_hd__a21oi_1 _10908_ (.A1(\CPU_Xreg_value_a4[14][24] ),
    .A2(_04697_),
    .B1(net91),
    .Y(_04959_));
 sky130_fd_sc_hd__a22oi_1 _10909_ (.A1(\CPU_Xreg_value_a4[10][24] ),
    .A2(_04733_),
    .B1(net18),
    .B2(\CPU_Xreg_value_a4[3][24] ),
    .Y(_04960_));
 sky130_fd_sc_hd__a22oi_1 _10910_ (.A1(\CPU_Xreg_value_a4[13][24] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][24] ),
    .Y(_04961_));
 sky130_fd_sc_hd__a22oi_1 _10911_ (.A1(\CPU_Xreg_value_a4[11][24] ),
    .A2(_04705_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][24] ),
    .Y(_04962_));
 sky130_fd_sc_hd__nand4_2 _10912_ (.A(_04959_),
    .B(_04960_),
    .C(_04961_),
    .D(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__a22o_1 _10913_ (.A1(\CPU_Xreg_value_a4[2][24] ),
    .A2(net22),
    .B1(net16),
    .B2(\CPU_Xreg_value_a4[1][24] ),
    .X(_04964_));
 sky130_fd_sc_hd__a221oi_1 _10914_ (.A1(\CPU_Xreg_value_a4[7][24] ),
    .A2(_04719_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][24] ),
    .C1(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__a22oi_1 _10915_ (.A1(\CPU_Xreg_value_a4[12][24] ),
    .A2(net26),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][24] ),
    .Y(_04966_));
 sky130_fd_sc_hd__a22oi_1 _10916_ (.A1(\CPU_Xreg_value_a4[15][24] ),
    .A2(_04729_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][24] ),
    .Y(_04967_));
 sky130_fd_sc_hd__nand3_1 _10917_ (.A(_04965_),
    .B(_04966_),
    .C(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__o22ai_4 _10918_ (.A1(net1542),
    .A2(_04692_),
    .B1(_04963_),
    .B2(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__mux2i_1 _10919_ (.A0(_04969_),
    .A1(_04511_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[24] ));
 sky130_fd_sc_hd__a21oi_1 _10920_ (.A1(net1696),
    .A2(_04729_),
    .B1(net91),
    .Y(_04970_));
 sky130_fd_sc_hd__a22oi_1 _10921_ (.A1(\CPU_Xreg_value_a4[14][25] ),
    .A2(_04697_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][25] ),
    .Y(_04971_));
 sky130_fd_sc_hd__a22oi_1 _10922_ (.A1(\CPU_Xreg_value_a4[7][25] ),
    .A2(_04719_),
    .B1(net26),
    .B2(net1692),
    .Y(_04972_));
 sky130_fd_sc_hd__a22oi_1 _10923_ (.A1(\CPU_Xreg_value_a4[10][25] ),
    .A2(_04733_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][25] ),
    .Y(_04973_));
 sky130_fd_sc_hd__nand4_1 _10924_ (.A(_04970_),
    .B(_04971_),
    .C(_04972_),
    .D(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__a22o_1 _10925_ (.A1(\CPU_Xreg_value_a4[2][25] ),
    .A2(net22),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][25] ),
    .X(_04975_));
 sky130_fd_sc_hd__a221oi_1 _10926_ (.A1(net1714),
    .A2(_04705_),
    .B1(net15),
    .B2(net1712),
    .C1(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__a22oi_1 _10927_ (.A1(\CPU_Xreg_value_a4[13][25] ),
    .A2(_04736_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][25] ),
    .Y(_04977_));
 sky130_fd_sc_hd__a22oi_1 _10928_ (.A1(net1719),
    .A2(net18),
    .B1(net16),
    .B2(net1695),
    .Y(_04978_));
 sky130_fd_sc_hd__nand3_1 _10929_ (.A(_04976_),
    .B(_04977_),
    .C(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__o22ai_1 _10930_ (.A1(net1279),
    .A2(_04692_),
    .B1(_04974_),
    .B2(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__mux2i_1 _10931_ (.A0(net1720),
    .A1(_04523_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[25] ));
 sky130_fd_sc_hd__a21oi_1 _10932_ (.A1(\CPU_Xreg_value_a4[9][26] ),
    .A2(_04711_),
    .B1(net90),
    .Y(_04981_));
 sky130_fd_sc_hd__a22oi_1 _10933_ (.A1(\CPU_Xreg_value_a4[3][26] ),
    .A2(net18),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][26] ),
    .Y(_04982_));
 sky130_fd_sc_hd__a22oi_1 _10934_ (.A1(\CPU_Xreg_value_a4[15][26] ),
    .A2(_04729_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][26] ),
    .Y(_04983_));
 sky130_fd_sc_hd__a22oi_1 _10935_ (.A1(\CPU_Xreg_value_a4[11][26] ),
    .A2(_04705_),
    .B1(net26),
    .B2(\CPU_Xreg_value_a4[12][26] ),
    .Y(_04984_));
 sky130_fd_sc_hd__nand4_1 _10936_ (.A(_04981_),
    .B(_04982_),
    .C(_04983_),
    .D(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__a22o_1 _10937_ (.A1(\CPU_Xreg_value_a4[10][26] ),
    .A2(_04733_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][26] ),
    .X(_04986_));
 sky130_fd_sc_hd__a221oi_1 _10938_ (.A1(\CPU_Xreg_value_a4[2][26] ),
    .A2(net22),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][26] ),
    .C1(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__a22oi_1 _10939_ (.A1(\CPU_Xreg_value_a4[1][26] ),
    .A2(net16),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][26] ),
    .Y(_04988_));
 sky130_fd_sc_hd__a22oi_1 _10940_ (.A1(\CPU_Xreg_value_a4[7][26] ),
    .A2(_04719_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][26] ),
    .Y(_04989_));
 sky130_fd_sc_hd__nand3_1 _10941_ (.A(_04987_),
    .B(_04988_),
    .C(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__o22ai_4 _10942_ (.A1(net1852),
    .A2(_04692_),
    .B1(_04985_),
    .B2(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_1 _10943_ (.A(_04535_),
    .B(_04752_),
    .Y(_04992_));
 sky130_fd_sc_hd__o21ai_0 _10944_ (.A1(_04752_),
    .A2(_04991_),
    .B1(_04992_),
    .Y(\CPU_src2_value_a2[26] ));
 sky130_fd_sc_hd__a21oi_1 _10945_ (.A1(\CPU_Xreg_value_a4[8][27] ),
    .A2(net24),
    .B1(net90),
    .Y(_04993_));
 sky130_fd_sc_hd__a22oi_1 _10946_ (.A1(\CPU_Xreg_value_a4[3][27] ),
    .A2(net19),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][27] ),
    .Y(_04994_));
 sky130_fd_sc_hd__a22oi_1 _10947_ (.A1(\CPU_Xreg_value_a4[2][27] ),
    .A2(net21),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][27] ),
    .Y(_04995_));
 sky130_fd_sc_hd__a22oi_1 _10948_ (.A1(\CPU_Xreg_value_a4[10][27] ),
    .A2(_04733_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][27] ),
    .Y(_04996_));
 sky130_fd_sc_hd__nand4_2 _10949_ (.A(_04993_),
    .B(_04994_),
    .C(_04995_),
    .D(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a22o_1 _10950_ (.A1(\CPU_Xreg_value_a4[1][27] ),
    .A2(net16),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][27] ),
    .X(_04998_));
 sky130_fd_sc_hd__a221oi_1 _10951_ (.A1(\CPU_Xreg_value_a4[7][27] ),
    .A2(_04719_),
    .B1(net25),
    .B2(\CPU_Xreg_value_a4[12][27] ),
    .C1(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__a22oi_1 _10952_ (.A1(\CPU_Xreg_value_a4[11][27] ),
    .A2(_04705_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][27] ),
    .Y(_05000_));
 sky130_fd_sc_hd__a22oi_1 _10953_ (.A1(\CPU_Xreg_value_a4[15][27] ),
    .A2(_04729_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][27] ),
    .Y(_05001_));
 sky130_fd_sc_hd__nand3_1 _10954_ (.A(_04999_),
    .B(_05000_),
    .C(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__o22ai_4 _10955_ (.A1(net1669),
    .A2(_04692_),
    .B1(_04997_),
    .B2(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__mux2i_1 _10956_ (.A0(_05003_),
    .A1(_03074_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[27] ));
 sky130_fd_sc_hd__a21oi_1 _10957_ (.A1(\CPU_Xreg_value_a4[1][28] ),
    .A2(net16),
    .B1(net91),
    .Y(_05004_));
 sky130_fd_sc_hd__a22oi_1 _10958_ (.A1(\CPU_Xreg_value_a4[6][28] ),
    .A2(_04740_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][28] ),
    .Y(_05005_));
 sky130_fd_sc_hd__a22oi_1 _10959_ (.A1(\CPU_Xreg_value_a4[7][28] ),
    .A2(_04719_),
    .B1(net26),
    .B2(\CPU_Xreg_value_a4[12][28] ),
    .Y(_05006_));
 sky130_fd_sc_hd__a22oi_1 _10960_ (.A1(\CPU_Xreg_value_a4[11][28] ),
    .A2(_04705_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][28] ),
    .Y(_05007_));
 sky130_fd_sc_hd__nand4_1 _10961_ (.A(_05004_),
    .B(_05005_),
    .C(_05006_),
    .D(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__a22o_1 _10962_ (.A1(\CPU_Xreg_value_a4[5][28] ),
    .A2(_04730_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][28] ),
    .X(_05009_));
 sky130_fd_sc_hd__a221oi_1 _10963_ (.A1(\CPU_Xreg_value_a4[2][28] ),
    .A2(net20),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][28] ),
    .C1(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__a22oi_1 _10964_ (.A1(\CPU_Xreg_value_a4[3][28] ),
    .A2(net18),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][28] ),
    .Y(_05011_));
 sky130_fd_sc_hd__a22oi_1 _10965_ (.A1(\CPU_Xreg_value_a4[10][28] ),
    .A2(_04733_),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][28] ),
    .Y(_05012_));
 sky130_fd_sc_hd__nand3_1 _10966_ (.A(_05010_),
    .B(_05011_),
    .C(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__o22ai_2 _10967_ (.A1(net1455),
    .A2(_04692_),
    .B1(_05008_),
    .B2(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__mux2i_1 _10968_ (.A0(_05014_),
    .A1(_03098_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[28] ));
 sky130_fd_sc_hd__a21oi_1 _10969_ (.A1(\CPU_Xreg_value_a4[4][29] ),
    .A2(_04742_),
    .B1(net91),
    .Y(_05015_));
 sky130_fd_sc_hd__a22oi_1 _10970_ (.A1(\CPU_Xreg_value_a4[15][29] ),
    .A2(_04729_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][29] ),
    .Y(_05016_));
 sky130_fd_sc_hd__a22oi_1 _10971_ (.A1(\CPU_Xreg_value_a4[12][29] ),
    .A2(net26),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][29] ),
    .Y(_05017_));
 sky130_fd_sc_hd__a22oi_1 _10972_ (.A1(\CPU_Xreg_value_a4[10][29] ),
    .A2(_04733_),
    .B1(net18),
    .B2(\CPU_Xreg_value_a4[3][29] ),
    .Y(_05018_));
 sky130_fd_sc_hd__nand4_1 _10973_ (.A(_05015_),
    .B(_05016_),
    .C(_05017_),
    .D(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__a22o_1 _10974_ (.A1(\CPU_Xreg_value_a4[1][29] ),
    .A2(net16),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][29] ),
    .X(_05020_));
 sky130_fd_sc_hd__a221oi_1 _10975_ (.A1(\CPU_Xreg_value_a4[11][29] ),
    .A2(_04705_),
    .B1(net22),
    .B2(\CPU_Xreg_value_a4[2][29] ),
    .C1(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__a22oi_1 _10976_ (.A1(\CPU_Xreg_value_a4[7][29] ),
    .A2(_04719_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][29] ),
    .Y(_05022_));
 sky130_fd_sc_hd__a22oi_1 _10977_ (.A1(\CPU_Xreg_value_a4[9][29] ),
    .A2(_04711_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][29] ),
    .Y(_05023_));
 sky130_fd_sc_hd__nand3_1 _10978_ (.A(_05021_),
    .B(_05022_),
    .C(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__o22ai_1 _10979_ (.A1(net1266),
    .A2(_04692_),
    .B1(_05019_),
    .B2(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_1 _10980_ (.A(_04752_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__a21o_1 _10981_ (.A1(_04559_),
    .A2(_04752_),
    .B1(_05026_),
    .X(\CPU_src2_value_a2[29] ));
 sky130_fd_sc_hd__a21oi_1 _10982_ (.A1(\CPU_Xreg_value_a4[14][2] ),
    .A2(_04697_),
    .B1(net90),
    .Y(_05027_));
 sky130_fd_sc_hd__a22oi_1 _10983_ (.A1(\CPU_Xreg_value_a4[2][2] ),
    .A2(net21),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][2] ),
    .Y(_05028_));
 sky130_fd_sc_hd__a22oi_1 _10984_ (.A1(\CPU_Xreg_value_a4[3][2] ),
    .A2(_04724_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][2] ),
    .Y(_05029_));
 sky130_fd_sc_hd__a22oi_1 _10985_ (.A1(\CPU_Xreg_value_a4[7][2] ),
    .A2(_04719_),
    .B1(_04707_),
    .B2(\CPU_Xreg_value_a4[12][2] ),
    .Y(_05030_));
 sky130_fd_sc_hd__nand4_2 _10986_ (.A(_05027_),
    .B(_05028_),
    .C(_05029_),
    .D(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__a22o_1 _10987_ (.A1(\CPU_Xreg_value_a4[13][2] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][2] ),
    .X(_05032_));
 sky130_fd_sc_hd__a221oi_1 _10988_ (.A1(\CPU_Xreg_value_a4[11][2] ),
    .A2(_04705_),
    .B1(_04726_),
    .B2(\CPU_Xreg_value_a4[1][2] ),
    .C1(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__a22oi_1 _10989_ (.A1(\CPU_Xreg_value_a4[15][2] ),
    .A2(_04729_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][2] ),
    .Y(_05034_));
 sky130_fd_sc_hd__a22oi_1 _10990_ (.A1(\CPU_Xreg_value_a4[8][2] ),
    .A2(_04713_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][2] ),
    .Y(_05035_));
 sky130_fd_sc_hd__nand3_1 _10991_ (.A(_05033_),
    .B(_05034_),
    .C(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__o22ai_4 _10992_ (.A1(net1666),
    .A2(_04692_),
    .B1(_05031_),
    .B2(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(\CPU_result_a3[2] ),
    .B(_04752_),
    .Y(_05038_));
 sky130_fd_sc_hd__o21ai_0 _10994_ (.A1(_04752_),
    .A2(_05037_),
    .B1(_05038_),
    .Y(\CPU_src2_value_a2[2] ));
 sky130_fd_sc_hd__a21oi_1 _10995_ (.A1(\CPU_Xreg_value_a4[9][30] ),
    .A2(_04711_),
    .B1(net91),
    .Y(_05039_));
 sky130_fd_sc_hd__a22oi_1 _10996_ (.A1(\CPU_Xreg_value_a4[2][30] ),
    .A2(net20),
    .B1(net15),
    .B2(\CPU_Xreg_value_a4[4][30] ),
    .Y(_05040_));
 sky130_fd_sc_hd__a22oi_1 _10997_ (.A1(\CPU_Xreg_value_a4[11][30] ),
    .A2(_04705_),
    .B1(_04719_),
    .B2(\CPU_Xreg_value_a4[7][30] ),
    .Y(_05041_));
 sky130_fd_sc_hd__a22oi_1 _10998_ (.A1(\CPU_Xreg_value_a4[3][30] ),
    .A2(net18),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][30] ),
    .Y(_05042_));
 sky130_fd_sc_hd__nand4_1 _10999_ (.A(_05039_),
    .B(_05040_),
    .C(_05041_),
    .D(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__a22o_1 _11000_ (.A1(\CPU_Xreg_value_a4[1][30] ),
    .A2(net16),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][30] ),
    .X(_05044_));
 sky130_fd_sc_hd__a221oi_1 _11001_ (.A1(\CPU_Xreg_value_a4[12][30] ),
    .A2(net25),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][30] ),
    .C1(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a22oi_1 _11002_ (.A1(\CPU_Xreg_value_a4[13][30] ),
    .A2(_04736_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][30] ),
    .Y(_05046_));
 sky130_fd_sc_hd__a22oi_1 _11003_ (.A1(\CPU_Xreg_value_a4[10][30] ),
    .A2(_04733_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][30] ),
    .Y(_05047_));
 sky130_fd_sc_hd__nand3_1 _11004_ (.A(_05045_),
    .B(_05046_),
    .C(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__o22ai_4 _11005_ (.A1(net1853),
    .A2(_04692_),
    .B1(_05043_),
    .B2(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__mux2i_1 _11006_ (.A0(_05049_),
    .A1(_03161_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[30] ));
 sky130_fd_sc_hd__a21oi_1 _11007_ (.A1(\CPU_Xreg_value_a4[8][31] ),
    .A2(net23),
    .B1(net92),
    .Y(_05050_));
 sky130_fd_sc_hd__a22oi_1 _11008_ (.A1(\CPU_Xreg_value_a4[7][31] ),
    .A2(_04719_),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][31] ),
    .Y(_05051_));
 sky130_fd_sc_hd__a22oi_1 _11009_ (.A1(\CPU_Xreg_value_a4[15][31] ),
    .A2(_04729_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][31] ),
    .Y(_05052_));
 sky130_fd_sc_hd__a22oi_1 _11010_ (.A1(\CPU_Xreg_value_a4[12][31] ),
    .A2(net25),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][31] ),
    .Y(_05053_));
 sky130_fd_sc_hd__nand4_1 _11011_ (.A(_05050_),
    .B(_05051_),
    .C(_05052_),
    .D(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__a22o_1 _11012_ (.A1(\CPU_Xreg_value_a4[1][31] ),
    .A2(net17),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][31] ),
    .X(_05055_));
 sky130_fd_sc_hd__a221oi_1 _11013_ (.A1(\CPU_Xreg_value_a4[2][31] ),
    .A2(net20),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][31] ),
    .C1(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__a22oi_1 _11014_ (.A1(\CPU_Xreg_value_a4[11][31] ),
    .A2(_04705_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][31] ),
    .Y(_05057_));
 sky130_fd_sc_hd__a22oi_1 _11015_ (.A1(\CPU_Xreg_value_a4[3][31] ),
    .A2(net19),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][31] ),
    .Y(_05058_));
 sky130_fd_sc_hd__nand3_1 _11016_ (.A(_05056_),
    .B(_05057_),
    .C(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__o22ai_4 _11017_ (.A1(net1683),
    .A2(_04692_),
    .B1(_05054_),
    .B2(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__mux2i_1 _11018_ (.A0(_05060_),
    .A1(_03189_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[31] ));
 sky130_fd_sc_hd__a21oi_1 _11019_ (.A1(\CPU_Xreg_value_a4[4][3] ),
    .A2(net14),
    .B1(net92),
    .Y(_05061_));
 sky130_fd_sc_hd__a22oi_1 _11020_ (.A1(\CPU_Xreg_value_a4[13][3] ),
    .A2(_04736_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][3] ),
    .Y(_05062_));
 sky130_fd_sc_hd__a22oi_1 _11021_ (.A1(\CPU_Xreg_value_a4[11][3] ),
    .A2(_04705_),
    .B1(_04724_),
    .B2(\CPU_Xreg_value_a4[3][3] ),
    .Y(_05063_));
 sky130_fd_sc_hd__a22oi_1 _11022_ (.A1(\CPU_Xreg_value_a4[15][3] ),
    .A2(_04729_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][3] ),
    .Y(_05064_));
 sky130_fd_sc_hd__nand4_2 _11023_ (.A(_05061_),
    .B(_05062_),
    .C(_05063_),
    .D(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__a22o_1 _11024_ (.A1(\CPU_Xreg_value_a4[2][3] ),
    .A2(_04716_),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][3] ),
    .X(_05066_));
 sky130_fd_sc_hd__a221oi_1 _11025_ (.A1(\CPU_Xreg_value_a4[7][3] ),
    .A2(_04719_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][3] ),
    .C1(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__a22oi_1 _11026_ (.A1(\CPU_Xreg_value_a4[9][3] ),
    .A2(_04711_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][3] ),
    .Y(_05068_));
 sky130_fd_sc_hd__a22oi_1 _11027_ (.A1(\CPU_Xreg_value_a4[12][3] ),
    .A2(_04707_),
    .B1(_04726_),
    .B2(\CPU_Xreg_value_a4[1][3] ),
    .Y(_05069_));
 sky130_fd_sc_hd__nand3_1 _11028_ (.A(_05067_),
    .B(_05068_),
    .C(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__o22ai_4 _11029_ (.A1(net1520),
    .A2(_04692_),
    .B1(_05065_),
    .B2(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(\CPU_result_a3[3] ),
    .B(_04752_),
    .Y(_05072_));
 sky130_fd_sc_hd__o21ai_0 _11031_ (.A1(_04752_),
    .A2(_05071_),
    .B1(_05072_),
    .Y(\CPU_src2_value_a2[3] ));
 sky130_fd_sc_hd__a21oi_1 _11032_ (.A1(\CPU_Xreg_value_a4[5][4] ),
    .A2(_04730_),
    .B1(net90),
    .Y(_05073_));
 sky130_fd_sc_hd__a22oi_1 _11033_ (.A1(\CPU_Xreg_value_a4[13][4] ),
    .A2(_04736_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][4] ),
    .Y(_05074_));
 sky130_fd_sc_hd__a22oi_1 _11034_ (.A1(\CPU_Xreg_value_a4[12][4] ),
    .A2(_04707_),
    .B1(_04724_),
    .B2(\CPU_Xreg_value_a4[3][4] ),
    .Y(_05075_));
 sky130_fd_sc_hd__a22oi_1 _11035_ (.A1(\CPU_Xreg_value_a4[10][4] ),
    .A2(_04733_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][4] ),
    .Y(_05076_));
 sky130_fd_sc_hd__nand4_2 _11036_ (.A(_05073_),
    .B(_05074_),
    .C(_05075_),
    .D(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__a22o_1 _11037_ (.A1(\CPU_Xreg_value_a4[7][4] ),
    .A2(_04719_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][4] ),
    .X(_05078_));
 sky130_fd_sc_hd__a221oi_1 _11038_ (.A1(\CPU_Xreg_value_a4[2][4] ),
    .A2(net21),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][4] ),
    .C1(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__a22oi_1 _11039_ (.A1(\CPU_Xreg_value_a4[11][4] ),
    .A2(_04705_),
    .B1(net24),
    .B2(\CPU_Xreg_value_a4[8][4] ),
    .Y(_05080_));
 sky130_fd_sc_hd__a22oi_1 _11040_ (.A1(\CPU_Xreg_value_a4[1][4] ),
    .A2(_04726_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][4] ),
    .Y(_05081_));
 sky130_fd_sc_hd__nand3_1 _11041_ (.A(_05079_),
    .B(_05080_),
    .C(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__o22ai_4 _11042_ (.A1(net1673),
    .A2(_04692_),
    .B1(_05077_),
    .B2(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _11043_ (.A(\CPU_result_a3[4] ),
    .B(_04752_),
    .Y(_05084_));
 sky130_fd_sc_hd__o21ai_0 _11044_ (.A1(_04752_),
    .A2(_05083_),
    .B1(_05084_),
    .Y(\CPU_src2_value_a2[4] ));
 sky130_fd_sc_hd__a21oi_1 _11045_ (.A1(\CPU_Xreg_value_a4[6][5] ),
    .A2(_04740_),
    .B1(net92),
    .Y(_05085_));
 sky130_fd_sc_hd__a22oi_1 _11046_ (.A1(\CPU_Xreg_value_a4[1][5] ),
    .A2(_04726_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][5] ),
    .Y(_05086_));
 sky130_fd_sc_hd__a22oi_1 _11047_ (.A1(\CPU_Xreg_value_a4[11][5] ),
    .A2(_04705_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][5] ),
    .Y(_05087_));
 sky130_fd_sc_hd__a22oi_1 _11048_ (.A1(\CPU_Xreg_value_a4[7][5] ),
    .A2(_04719_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][5] ),
    .Y(_05088_));
 sky130_fd_sc_hd__nand4_2 _11049_ (.A(_05085_),
    .B(_05086_),
    .C(_05087_),
    .D(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a22o_1 _11050_ (.A1(\CPU_Xreg_value_a4[9][5] ),
    .A2(_04711_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][5] ),
    .X(_05090_));
 sky130_fd_sc_hd__a221oi_1 _11051_ (.A1(\CPU_Xreg_value_a4[2][5] ),
    .A2(net21),
    .B1(_04733_),
    .B2(\CPU_Xreg_value_a4[10][5] ),
    .C1(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a22oi_1 _11052_ (.A1(\CPU_Xreg_value_a4[3][5] ),
    .A2(net19),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][5] ),
    .Y(_05092_));
 sky130_fd_sc_hd__a22oi_1 _11053_ (.A1(\CPU_Xreg_value_a4[12][5] ),
    .A2(net25),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][5] ),
    .Y(_05093_));
 sky130_fd_sc_hd__nand3_1 _11054_ (.A(_05091_),
    .B(_05092_),
    .C(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__o22ai_4 _11055_ (.A1(net1618),
    .A2(_04692_),
    .B1(_05089_),
    .B2(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__mux2i_1 _11056_ (.A0(_05095_),
    .A1(_03217_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[5] ));
 sky130_fd_sc_hd__a21oi_1 _11057_ (.A1(\CPU_Xreg_value_a4[4][6] ),
    .A2(net14),
    .B1(net90),
    .Y(_05096_));
 sky130_fd_sc_hd__a22oi_1 _11058_ (.A1(\CPU_Xreg_value_a4[12][6] ),
    .A2(net25),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][6] ),
    .Y(_05097_));
 sky130_fd_sc_hd__a22oi_1 _11059_ (.A1(\CPU_Xreg_value_a4[3][6] ),
    .A2(net19),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][6] ),
    .Y(_05098_));
 sky130_fd_sc_hd__a22oi_1 _11060_ (.A1(\CPU_Xreg_value_a4[11][6] ),
    .A2(_04705_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][6] ),
    .Y(_05099_));
 sky130_fd_sc_hd__nand4_2 _11061_ (.A(_05096_),
    .B(_05097_),
    .C(_05098_),
    .D(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__a22o_1 _11062_ (.A1(\CPU_Xreg_value_a4[10][6] ),
    .A2(_04733_),
    .B1(net23),
    .B2(\CPU_Xreg_value_a4[8][6] ),
    .X(_05101_));
 sky130_fd_sc_hd__a221oi_1 _11063_ (.A1(\CPU_Xreg_value_a4[7][6] ),
    .A2(_04719_),
    .B1(net16),
    .B2(\CPU_Xreg_value_a4[1][6] ),
    .C1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__a22oi_1 _11064_ (.A1(\CPU_Xreg_value_a4[2][6] ),
    .A2(net21),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][6] ),
    .Y(_05103_));
 sky130_fd_sc_hd__a22oi_1 _11065_ (.A1(\CPU_Xreg_value_a4[6][6] ),
    .A2(_04740_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][6] ),
    .Y(_05104_));
 sky130_fd_sc_hd__nand3_1 _11066_ (.A(_05102_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__o22ai_4 _11067_ (.A1(\CPU_Xreg_value_a4[0][6] ),
    .A2(_04692_),
    .B1(_05100_),
    .B2(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__mux2i_1 _11068_ (.A0(_05106_),
    .A1(_03225_),
    .S(_04752_),
    .Y(\CPU_src2_value_a2[6] ));
 sky130_fd_sc_hd__a21oi_1 _11069_ (.A1(\CPU_Xreg_value_a4[10][7] ),
    .A2(_04733_),
    .B1(net92),
    .Y(_05107_));
 sky130_fd_sc_hd__a22oi_1 _11070_ (.A1(\CPU_Xreg_value_a4[7][7] ),
    .A2(_04719_),
    .B1(_04729_),
    .B2(\CPU_Xreg_value_a4[15][7] ),
    .Y(_05108_));
 sky130_fd_sc_hd__a22oi_1 _11071_ (.A1(\CPU_Xreg_value_a4[12][7] ),
    .A2(_04707_),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][7] ),
    .Y(_05109_));
 sky130_fd_sc_hd__a22oi_1 _11072_ (.A1(\CPU_Xreg_value_a4[14][7] ),
    .A2(_04697_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][7] ),
    .Y(_05110_));
 sky130_fd_sc_hd__nand4_1 _11073_ (.A(_05107_),
    .B(_05108_),
    .C(_05109_),
    .D(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__a22o_1 _11074_ (.A1(\CPU_Xreg_value_a4[1][7] ),
    .A2(_04726_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][7] ),
    .X(_05112_));
 sky130_fd_sc_hd__a221oi_1 _11075_ (.A1(\CPU_Xreg_value_a4[2][7] ),
    .A2(_04716_),
    .B1(_04724_),
    .B2(\CPU_Xreg_value_a4[3][7] ),
    .C1(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__a22oi_1 _11076_ (.A1(\CPU_Xreg_value_a4[13][7] ),
    .A2(_04736_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][7] ),
    .Y(_05114_));
 sky130_fd_sc_hd__a22oi_1 _11077_ (.A1(\CPU_Xreg_value_a4[11][7] ),
    .A2(_04705_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][7] ),
    .Y(_05115_));
 sky130_fd_sc_hd__nand3_1 _11078_ (.A(_05113_),
    .B(_05114_),
    .C(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__o22ai_4 _11079_ (.A1(\CPU_Xreg_value_a4[0][7] ),
    .A2(_04692_),
    .B1(_05111_),
    .B2(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(_03235_),
    .B(_04752_),
    .Y(_05118_));
 sky130_fd_sc_hd__o21ai_0 _11081_ (.A1(_04752_),
    .A2(_05117_),
    .B1(_05118_),
    .Y(\CPU_src2_value_a2[7] ));
 sky130_fd_sc_hd__a21oi_1 _11082_ (.A1(\CPU_Xreg_value_a4[3][8] ),
    .A2(net19),
    .B1(net90),
    .Y(_05119_));
 sky130_fd_sc_hd__a22oi_1 _11083_ (.A1(\CPU_Xreg_value_a4[11][8] ),
    .A2(_04705_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][8] ),
    .Y(_05120_));
 sky130_fd_sc_hd__a22oi_1 _11084_ (.A1(\CPU_Xreg_value_a4[1][8] ),
    .A2(_04726_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][8] ),
    .Y(_05121_));
 sky130_fd_sc_hd__a22oi_1 _11085_ (.A1(\CPU_Xreg_value_a4[6][8] ),
    .A2(_04740_),
    .B1(_04730_),
    .B2(\CPU_Xreg_value_a4[5][8] ),
    .Y(_05122_));
 sky130_fd_sc_hd__nand4_1 _11086_ (.A(_05119_),
    .B(_05120_),
    .C(_05121_),
    .D(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__a22o_1 _11087_ (.A1(\CPU_Xreg_value_a4[15][8] ),
    .A2(_04729_),
    .B1(_04736_),
    .B2(\CPU_Xreg_value_a4[13][8] ),
    .X(_05124_));
 sky130_fd_sc_hd__a221oi_1 _11088_ (.A1(\CPU_Xreg_value_a4[2][8] ),
    .A2(net21),
    .B1(_04719_),
    .B2(\CPU_Xreg_value_a4[7][8] ),
    .C1(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__a22oi_1 _11089_ (.A1(\CPU_Xreg_value_a4[10][8] ),
    .A2(_04733_),
    .B1(net14),
    .B2(\CPU_Xreg_value_a4[4][8] ),
    .Y(_05126_));
 sky130_fd_sc_hd__a22oi_1 _11090_ (.A1(\CPU_Xreg_value_a4[12][8] ),
    .A2(net25),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][8] ),
    .Y(_05127_));
 sky130_fd_sc_hd__nand3_1 _11091_ (.A(_05125_),
    .B(_05126_),
    .C(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__o22ai_4 _11092_ (.A1(net1674),
    .A2(_04692_),
    .B1(_05123_),
    .B2(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _11093_ (.A(_03248_),
    .B(_04752_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_0 _11094_ (.A1(_04752_),
    .A2(_05129_),
    .B1(_05130_),
    .Y(\CPU_src2_value_a2[8] ));
 sky130_fd_sc_hd__a21oi_1 _11095_ (.A1(\CPU_Xreg_value_a4[5][9] ),
    .A2(_04730_),
    .B1(net92),
    .Y(_05131_));
 sky130_fd_sc_hd__a22oi_1 _11096_ (.A1(\CPU_Xreg_value_a4[13][9] ),
    .A2(_04736_),
    .B1(_04713_),
    .B2(\CPU_Xreg_value_a4[8][9] ),
    .Y(_05132_));
 sky130_fd_sc_hd__a22oi_1 _11097_ (.A1(\CPU_Xreg_value_a4[15][9] ),
    .A2(_04729_),
    .B1(_04711_),
    .B2(\CPU_Xreg_value_a4[9][9] ),
    .Y(_05133_));
 sky130_fd_sc_hd__a22oi_1 _11098_ (.A1(\CPU_Xreg_value_a4[11][9] ),
    .A2(_04705_),
    .B1(_04742_),
    .B2(\CPU_Xreg_value_a4[4][9] ),
    .Y(_05134_));
 sky130_fd_sc_hd__nand4_2 _11099_ (.A(_05131_),
    .B(_05132_),
    .C(_05133_),
    .D(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__a22o_1 _11100_ (.A1(\CPU_Xreg_value_a4[10][9] ),
    .A2(_04733_),
    .B1(_04726_),
    .B2(\CPU_Xreg_value_a4[1][9] ),
    .X(_05136_));
 sky130_fd_sc_hd__a221oi_1 _11101_ (.A1(\CPU_Xreg_value_a4[2][9] ),
    .A2(_04716_),
    .B1(_04697_),
    .B2(\CPU_Xreg_value_a4[14][9] ),
    .C1(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__a22oi_1 _11102_ (.A1(\CPU_Xreg_value_a4[7][9] ),
    .A2(_04719_),
    .B1(net25),
    .B2(\CPU_Xreg_value_a4[12][9] ),
    .Y(_05138_));
 sky130_fd_sc_hd__a22oi_1 _11103_ (.A1(\CPU_Xreg_value_a4[3][9] ),
    .A2(_04724_),
    .B1(_04740_),
    .B2(\CPU_Xreg_value_a4[6][9] ),
    .Y(_05139_));
 sky130_fd_sc_hd__nand3_1 _11104_ (.A(_05137_),
    .B(_05138_),
    .C(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__o22ai_4 _11105_ (.A1(net1678),
    .A2(_04692_),
    .B1(_05135_),
    .B2(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(_03258_),
    .B(_04752_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_0 _11107_ (.A1(_04752_),
    .A2(_05141_),
    .B1(_05142_),
    .Y(\CPU_src2_value_a2[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__a21oi_1 _11111_ (.A1(net1139),
    .A2(_02400_),
    .B1(net101),
    .Y(_05146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__a22oi_1 _11114_ (.A1(net1251),
    .A2(_01553_),
    .B1(_02247_),
    .B2(net1237),
    .Y(_05149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__a22oi_1 _11117_ (.A1(net551),
    .A2(net80),
    .B1(net73),
    .B2(net1114),
    .Y(_05152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__a22oi_1 _11120_ (.A1(net519),
    .A2(_01631_),
    .B1(net65),
    .B2(net715),
    .Y(_05155_));
 sky130_fd_sc_hd__nand4_1 _11121_ (.A(_05146_),
    .B(_05149_),
    .C(_05152_),
    .D(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__a22oi_1 _11124_ (.A1(net785),
    .A2(_01322_),
    .B1(_02092_),
    .B2(net1313),
    .Y(_05159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__a22oi_1 _11127_ (.A1(net1413),
    .A2(net63),
    .B1(net44),
    .B2(net401),
    .Y(_05162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__a22oi_1 _11131_ (.A1(net1204),
    .A2(_01705_),
    .B1(net54),
    .B2(net1050),
    .Y(_05166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__a22oi_1 _11134_ (.A1(net980),
    .A2(_01397_),
    .B1(_02172_),
    .B2(net650),
    .Y(_05169_));
 sky130_fd_sc_hd__nand4_1 _11135_ (.A(_05159_),
    .B(_05162_),
    .C(_05166_),
    .D(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__o22a_1 _11136_ (.A1(net848),
    .A2(_01170_),
    .B1(_05156_),
    .B2(_05170_),
    .X(\w_CPU_dmem_rd_data_a4[0] ));
 sky130_fd_sc_hd__a21oi_1 _11137_ (.A1(net1195),
    .A2(_02400_),
    .B1(net99),
    .Y(_05171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__a22oi_1 _11139_ (.A1(net456),
    .A2(_01322_),
    .B1(net43),
    .B2(net990),
    .Y(_05173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__a22oi_1 _11142_ (.A1(net1129),
    .A2(_01553_),
    .B1(_02092_),
    .B2(net1310),
    .Y(_05176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__a22oi_1 _11145_ (.A1(net393),
    .A2(_01397_),
    .B1(net81),
    .B2(net437),
    .Y(_05179_));
 sky130_fd_sc_hd__nand4_1 _11146_ (.A(_05171_),
    .B(_05173_),
    .C(_05176_),
    .D(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__a22o_1 _11148_ (.A1(net966),
    .A2(net55),
    .B1(_02247_),
    .B2(net666),
    .X(_05182_));
 sky130_fd_sc_hd__a221oi_1 _11149_ (.A1(net351),
    .A2(_01631_),
    .B1(net64),
    .B2(net924),
    .C1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__a22oi_1 _11151_ (.A1(net731),
    .A2(_01705_),
    .B1(net62),
    .B2(net273),
    .Y(_05185_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__a22oi_1 _11153_ (.A1(net612),
    .A2(net72),
    .B1(_02172_),
    .B2(net339),
    .Y(_05187_));
 sky130_fd_sc_hd__nand3_1 _11154_ (.A(_05183_),
    .B(_05185_),
    .C(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__o22a_1 _11155_ (.A1(net500),
    .A2(_01170_),
    .B1(_05180_),
    .B2(_05188_),
    .X(\w_CPU_dmem_rd_data_a4[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__a21oi_1 _11157_ (.A1(net323),
    .A2(_02247_),
    .B1(net99),
    .Y(_05190_));
 sky130_fd_sc_hd__a22oi_1 _11158_ (.A1(\CPU_Dmem_value_a5[12][11] ),
    .A2(net81),
    .B1(net72),
    .B2(\CPU_Dmem_value_a5[1][11] ),
    .Y(_05191_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__a22oi_1 _11160_ (.A1(\CPU_Dmem_value_a5[15][11] ),
    .A2(_01705_),
    .B1(net43),
    .B2(\CPU_Dmem_value_a5[8][11] ),
    .Y(_05193_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__a22oi_1 _11163_ (.A1(\CPU_Dmem_value_a5[10][11] ),
    .A2(_01322_),
    .B1(_01553_),
    .B2(\CPU_Dmem_value_a5[13][11] ),
    .Y(_05196_));
 sky130_fd_sc_hd__nand4_1 _11164_ (.A(_05190_),
    .B(_05191_),
    .C(_05193_),
    .D(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__a22o_1 _11166_ (.A1(\CPU_Dmem_value_a5[4][11] ),
    .A2(net55),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][11] ),
    .X(_05199_));
 sky130_fd_sc_hd__a221oi_1 _11167_ (.A1(net783),
    .A2(_01631_),
    .B1(net62),
    .B2(net381),
    .C1(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__a22oi_1 _11169_ (.A1(\CPU_Dmem_value_a5[11][11] ),
    .A2(_01397_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][11] ),
    .Y(_05202_));
 sky130_fd_sc_hd__a22oi_1 _11170_ (.A1(net1732),
    .A2(net64),
    .B1(_02172_),
    .B2(net225),
    .Y(_05203_));
 sky130_fd_sc_hd__nand3_1 _11171_ (.A(_05200_),
    .B(_05202_),
    .C(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__o22a_1 _11172_ (.A1(net299),
    .A2(_01170_),
    .B1(_05197_),
    .B2(_05204_),
    .X(\w_CPU_dmem_rd_data_a4[11] ));
 sky130_fd_sc_hd__a21oi_1 _11173_ (.A1(net840),
    .A2(_02247_),
    .B1(net100),
    .Y(_05205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__a22oi_1 _11175_ (.A1(\CPU_Dmem_value_a5[15][12] ),
    .A2(_01705_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][12] ),
    .Y(_05207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__a22oi_1 _11178_ (.A1(\CPU_Dmem_value_a5[11][12] ),
    .A2(_01397_),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][12] ),
    .Y(_05210_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__a22oi_1 _11181_ (.A1(\CPU_Dmem_value_a5[10][12] ),
    .A2(_01322_),
    .B1(_01631_),
    .B2(\CPU_Dmem_value_a5[14][12] ),
    .Y(_05213_));
 sky130_fd_sc_hd__nand4_1 _11182_ (.A(_05205_),
    .B(_05207_),
    .C(_05210_),
    .D(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__a22o_1 _11184_ (.A1(\CPU_Dmem_value_a5[3][12] ),
    .A2(net63),
    .B1(net54),
    .B2(\CPU_Dmem_value_a5[4][12] ),
    .X(_05216_));
 sky130_fd_sc_hd__a221oi_1 _11185_ (.A1(\CPU_Dmem_value_a5[1][12] ),
    .A2(net73),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][12] ),
    .C1(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__a22oi_1 _11187_ (.A1(\CPU_Dmem_value_a5[13][12] ),
    .A2(_01553_),
    .B1(net65),
    .B2(\CPU_Dmem_value_a5[2][12] ),
    .Y(_05219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__a22oi_1 _11189_ (.A1(\CPU_Dmem_value_a5[12][12] ),
    .A2(net80),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][12] ),
    .Y(_05221_));
 sky130_fd_sc_hd__nand3_1 _11190_ (.A(_05217_),
    .B(_05219_),
    .C(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__o22a_2 _11191_ (.A1(net371),
    .A2(_01170_),
    .B1(_05214_),
    .B2(_05222_),
    .X(\w_CPU_dmem_rd_data_a4[12] ));
 sky130_fd_sc_hd__a21oi_1 _11192_ (.A1(net1095),
    .A2(_02172_),
    .B1(net100),
    .Y(_05223_));
 sky130_fd_sc_hd__a22oi_1 _11193_ (.A1(\CPU_Dmem_value_a5[10][13] ),
    .A2(_01322_),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][13] ),
    .Y(_05224_));
 sky130_fd_sc_hd__a22oi_1 _11194_ (.A1(\CPU_Dmem_value_a5[15][13] ),
    .A2(_01705_),
    .B1(net64),
    .B2(\CPU_Dmem_value_a5[2][13] ),
    .Y(_05225_));
 sky130_fd_sc_hd__a22oi_1 _11195_ (.A1(\CPU_Dmem_value_a5[11][13] ),
    .A2(_01397_),
    .B1(_01631_),
    .B2(\CPU_Dmem_value_a5[14][13] ),
    .Y(_05226_));
 sky130_fd_sc_hd__nand4_1 _11196_ (.A(_05223_),
    .B(_05224_),
    .C(_05225_),
    .D(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__a22o_1 _11198_ (.A1(\CPU_Dmem_value_a5[3][13] ),
    .A2(net63),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][13] ),
    .X(_05229_));
 sky130_fd_sc_hd__a221oi_1 _11199_ (.A1(\CPU_Dmem_value_a5[12][13] ),
    .A2(net80),
    .B1(net73),
    .B2(\CPU_Dmem_value_a5[1][13] ),
    .C1(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__a22oi_1 _11200_ (.A1(\CPU_Dmem_value_a5[13][13] ),
    .A2(_01553_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][13] ),
    .Y(_05231_));
 sky130_fd_sc_hd__a22oi_1 _11201_ (.A1(\CPU_Dmem_value_a5[4][13] ),
    .A2(net54),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][13] ),
    .Y(_05232_));
 sky130_fd_sc_hd__nand3_1 _11202_ (.A(_05230_),
    .B(_05231_),
    .C(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__o22a_1 _11203_ (.A1(net537),
    .A2(_01170_),
    .B1(_05227_),
    .B2(_05233_),
    .X(\w_CPU_dmem_rd_data_a4[13] ));
 sky130_fd_sc_hd__a21oi_1 _11204_ (.A1(net219),
    .A2(_02400_),
    .B1(net99),
    .Y(_05234_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__a22oi_1 _11206_ (.A1(\CPU_Dmem_value_a5[14][14] ),
    .A2(_01631_),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][14] ),
    .Y(_05236_));
 sky130_fd_sc_hd__a22oi_1 _11207_ (.A1(\CPU_Dmem_value_a5[10][14] ),
    .A2(_01322_),
    .B1(net62),
    .B2(\CPU_Dmem_value_a5[3][14] ),
    .Y(_05237_));
 sky130_fd_sc_hd__a22oi_1 _11208_ (.A1(\CPU_Dmem_value_a5[11][14] ),
    .A2(_01397_),
    .B1(_01553_),
    .B2(\CPU_Dmem_value_a5[13][14] ),
    .Y(_05238_));
 sky130_fd_sc_hd__nand4_1 _11209_ (.A(_05234_),
    .B(_05236_),
    .C(_05237_),
    .D(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__a22o_1 _11210_ (.A1(\CPU_Dmem_value_a5[5][14] ),
    .A2(_02092_),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][14] ),
    .X(_05240_));
 sky130_fd_sc_hd__a221oi_1 _11211_ (.A1(\CPU_Dmem_value_a5[12][14] ),
    .A2(net80),
    .B1(net73),
    .B2(\CPU_Dmem_value_a5[1][14] ),
    .C1(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__a22oi_1 _11212_ (.A1(\CPU_Dmem_value_a5[15][14] ),
    .A2(_01705_),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][14] ),
    .Y(_05242_));
 sky130_fd_sc_hd__a22oi_1 _11213_ (.A1(\CPU_Dmem_value_a5[2][14] ),
    .A2(net65),
    .B1(net54),
    .B2(\CPU_Dmem_value_a5[4][14] ),
    .Y(_05243_));
 sky130_fd_sc_hd__nand3_1 _11214_ (.A(_05241_),
    .B(_05242_),
    .C(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__o22a_1 _11215_ (.A1(net315),
    .A2(_01170_),
    .B1(_05239_),
    .B2(_05244_),
    .X(\w_CPU_dmem_rd_data_a4[14] ));
 sky130_fd_sc_hd__a21oi_1 _11216_ (.A1(net421),
    .A2(_02172_),
    .B1(net99),
    .Y(_05245_));
 sky130_fd_sc_hd__a22oi_1 _11217_ (.A1(net694),
    .A2(_01553_),
    .B1(_01705_),
    .B2(net1028),
    .Y(_05246_));
 sky130_fd_sc_hd__a22oi_1 _11218_ (.A1(net952),
    .A2(_01322_),
    .B1(_02400_),
    .B2(net1048),
    .Y(_05247_));
 sky130_fd_sc_hd__a22oi_1 _11219_ (.A1(net515),
    .A2(_01631_),
    .B1(net72),
    .B2(net733),
    .Y(_05248_));
 sky130_fd_sc_hd__nand4_1 _11220_ (.A(_05245_),
    .B(_05246_),
    .C(_05247_),
    .D(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__a22o_1 _11221_ (.A1(\CPU_Dmem_value_a5[4][15] ),
    .A2(net55),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][15] ),
    .X(_05250_));
 sky130_fd_sc_hd__a221oi_1 _11222_ (.A1(net817),
    .A2(net64),
    .B1(net62),
    .B2(net825),
    .C1(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__a22oi_1 _11223_ (.A1(net1121),
    .A2(net80),
    .B1(_02092_),
    .B2(net353),
    .Y(_05252_));
 sky130_fd_sc_hd__a22oi_1 _11224_ (.A1(net632),
    .A2(_01397_),
    .B1(net43),
    .B2(net267),
    .Y(_05253_));
 sky130_fd_sc_hd__nand3_1 _11225_ (.A(_05251_),
    .B(_05252_),
    .C(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__o22a_1 _11226_ (.A1(net472),
    .A2(_01170_),
    .B1(_05249_),
    .B2(_05254_),
    .X(\w_CPU_dmem_rd_data_a4[15] ));
 sky130_fd_sc_hd__a21oi_1 _11227_ (.A1(net717),
    .A2(_02247_),
    .B1(net101),
    .Y(_05255_));
 sky130_fd_sc_hd__a22oi_1 _11228_ (.A1(net711),
    .A2(_01553_),
    .B1(net43),
    .B2(net1055),
    .Y(_05256_));
 sky130_fd_sc_hd__a22oi_1 _11229_ (.A1(net978),
    .A2(_01397_),
    .B1(net63),
    .B2(net998),
    .Y(_05257_));
 sky130_fd_sc_hd__a22oi_1 _11230_ (.A1(net942),
    .A2(_01322_),
    .B1(net65),
    .B2(net395),
    .Y(_05258_));
 sky130_fd_sc_hd__nand4_1 _11231_ (.A(_05255_),
    .B(_05256_),
    .C(_05257_),
    .D(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a22o_1 _11232_ (.A1(net709),
    .A2(_02092_),
    .B1(_02172_),
    .B2(net846),
    .X(_05260_));
 sky130_fd_sc_hd__a221oi_1 _11233_ (.A1(net801),
    .A2(net80),
    .B1(_01631_),
    .B2(net1087),
    .C1(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__a22oi_1 _11234_ (.A1(net391),
    .A2(net73),
    .B1(_02400_),
    .B2(net245),
    .Y(_05262_));
 sky130_fd_sc_hd__a22oi_1 _11235_ (.A1(net1210),
    .A2(_01705_),
    .B1(net55),
    .B2(net423),
    .Y(_05263_));
 sky130_fd_sc_hd__nand3_1 _11236_ (.A(_05261_),
    .B(_05262_),
    .C(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__o22a_1 _11237_ (.A1(net1162),
    .A2(_01170_),
    .B1(_05259_),
    .B2(_05264_),
    .X(\w_CPU_dmem_rd_data_a4[16] ));
 sky130_fd_sc_hd__a21oi_1 _11238_ (.A1(net1830),
    .A2(_02400_),
    .B1(net100),
    .Y(_05265_));
 sky130_fd_sc_hd__a22oi_1 _11239_ (.A1(\CPU_Dmem_value_a5[11][17] ),
    .A2(_01397_),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][17] ),
    .Y(_05266_));
 sky130_fd_sc_hd__a22oi_1 _11240_ (.A1(\CPU_Dmem_value_a5[14][17] ),
    .A2(_01631_),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][17] ),
    .Y(_05267_));
 sky130_fd_sc_hd__a22oi_1 _11241_ (.A1(\CPU_Dmem_value_a5[10][17] ),
    .A2(_01322_),
    .B1(net80),
    .B2(\CPU_Dmem_value_a5[12][17] ),
    .Y(_05268_));
 sky130_fd_sc_hd__nand4_1 _11242_ (.A(_05265_),
    .B(_05266_),
    .C(_05267_),
    .D(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a22o_1 _11243_ (.A1(\CPU_Dmem_value_a5[3][17] ),
    .A2(net63),
    .B1(net54),
    .B2(\CPU_Dmem_value_a5[4][17] ),
    .X(_05270_));
 sky130_fd_sc_hd__a221oi_1 _11244_ (.A1(\CPU_Dmem_value_a5[1][17] ),
    .A2(net73),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][17] ),
    .C1(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__a22oi_1 _11245_ (.A1(\CPU_Dmem_value_a5[13][17] ),
    .A2(_01553_),
    .B1(net65),
    .B2(\CPU_Dmem_value_a5[2][17] ),
    .Y(_05272_));
 sky130_fd_sc_hd__a22oi_1 _11246_ (.A1(\CPU_Dmem_value_a5[15][17] ),
    .A2(_01705_),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][17] ),
    .Y(_05273_));
 sky130_fd_sc_hd__nand3_1 _11247_ (.A(_05271_),
    .B(_05272_),
    .C(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__o22a_1 _11248_ (.A1(net741),
    .A2(_01170_),
    .B1(_05269_),
    .B2(_05274_),
    .X(\w_CPU_dmem_rd_data_a4[17] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__a21oi_1 _11250_ (.A1(net498),
    .A2(_02247_),
    .B1(net100),
    .Y(_05276_));
 sky130_fd_sc_hd__a22oi_1 _11251_ (.A1(\CPU_Dmem_value_a5[12][18] ),
    .A2(net80),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][18] ),
    .Y(_05277_));
 sky130_fd_sc_hd__a22oi_1 _11252_ (.A1(\CPU_Dmem_value_a5[11][18] ),
    .A2(_01397_),
    .B1(net64),
    .B2(\CPU_Dmem_value_a5[2][18] ),
    .Y(_05278_));
 sky130_fd_sc_hd__a22oi_1 _11253_ (.A1(\CPU_Dmem_value_a5[13][18] ),
    .A2(_01553_),
    .B1(_01705_),
    .B2(\CPU_Dmem_value_a5[15][18] ),
    .Y(_05279_));
 sky130_fd_sc_hd__nand4_1 _11254_ (.A(_05276_),
    .B(_05277_),
    .C(_05278_),
    .D(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__a22o_1 _11255_ (.A1(\CPU_Dmem_value_a5[1][18] ),
    .A2(net73),
    .B1(net63),
    .B2(\CPU_Dmem_value_a5[3][18] ),
    .X(_05281_));
 sky130_fd_sc_hd__a221oi_1 _11256_ (.A1(net1786),
    .A2(net54),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][18] ),
    .C1(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__a22oi_1 _11257_ (.A1(\CPU_Dmem_value_a5[10][18] ),
    .A2(_01322_),
    .B1(_02172_),
    .B2(net331),
    .Y(_05283_));
 sky130_fd_sc_hd__a22oi_1 _11258_ (.A1(\CPU_Dmem_value_a5[14][18] ),
    .A2(_01631_),
    .B1(_02400_),
    .B2(net567),
    .Y(_05284_));
 sky130_fd_sc_hd__nand3_1 _11259_ (.A(net1787),
    .B(_05283_),
    .C(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__o22a_2 _11260_ (.A1(net1018),
    .A2(_01170_),
    .B1(_05280_),
    .B2(net1788),
    .X(\w_CPU_dmem_rd_data_a4[18] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__a21oi_1 _11262_ (.A1(\CPU_Dmem_value_a5[7][19] ),
    .A2(_02247_),
    .B1(net100),
    .Y(_05287_));
 sky130_fd_sc_hd__a22oi_1 _11263_ (.A1(\CPU_Dmem_value_a5[13][19] ),
    .A2(_01553_),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][19] ),
    .Y(_05288_));
 sky130_fd_sc_hd__a22oi_1 _11264_ (.A1(\CPU_Dmem_value_a5[12][19] ),
    .A2(net81),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][19] ),
    .Y(_05289_));
 sky130_fd_sc_hd__a22oi_1 _11265_ (.A1(\CPU_Dmem_value_a5[10][19] ),
    .A2(_01322_),
    .B1(net62),
    .B2(\CPU_Dmem_value_a5[3][19] ),
    .Y(_05290_));
 sky130_fd_sc_hd__nand4_1 _11266_ (.A(_05287_),
    .B(_05288_),
    .C(_05289_),
    .D(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__a22oi_1 _11267_ (.A1(\CPU_Dmem_value_a5[11][19] ),
    .A2(_01397_),
    .B1(_02092_),
    .B2(net1036),
    .Y(_05292_));
 sky130_fd_sc_hd__a22oi_1 _11268_ (.A1(\CPU_Dmem_value_a5[2][19] ),
    .A2(net64),
    .B1(net54),
    .B2(\CPU_Dmem_value_a5[4][19] ),
    .Y(_05293_));
 sky130_fd_sc_hd__a22oi_1 _11269_ (.A1(\CPU_Dmem_value_a5[15][19] ),
    .A2(_01705_),
    .B1(net73),
    .B2(\CPU_Dmem_value_a5[1][19] ),
    .Y(_05294_));
 sky130_fd_sc_hd__a22oi_1 _11270_ (.A1(\CPU_Dmem_value_a5[14][19] ),
    .A2(_01631_),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][19] ),
    .Y(_05295_));
 sky130_fd_sc_hd__nand4_1 _11271_ (.A(_05292_),
    .B(_05293_),
    .C(_05294_),
    .D(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__o22a_2 _11272_ (.A1(net543),
    .A2(_01170_),
    .B1(_05291_),
    .B2(_05296_),
    .X(\w_CPU_dmem_rd_data_a4[19] ));
 sky130_fd_sc_hd__a21oi_1 _11273_ (.A1(net934),
    .A2(_02092_),
    .B1(net101),
    .Y(_05297_));
 sky130_fd_sc_hd__a22oi_1 _11274_ (.A1(net1208),
    .A2(_01397_),
    .B1(_01782_),
    .B2(net882),
    .Y(_05298_));
 sky130_fd_sc_hd__a22oi_1 _11275_ (.A1(net787),
    .A2(_01478_),
    .B1(_02018_),
    .B2(net271),
    .Y(_05299_));
 sky130_fd_sc_hd__a22oi_1 _11276_ (.A1(net1300),
    .A2(_01631_),
    .B1(_01861_),
    .B2(net1259),
    .Y(_05300_));
 sky130_fd_sc_hd__nand4_1 _11277_ (.A(_05297_),
    .B(_05298_),
    .C(_05299_),
    .D(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__a22o_1 _11278_ (.A1(\CPU_Dmem_value_a5[15][1] ),
    .A2(_01705_),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][1] ),
    .X(_05302_));
 sky130_fd_sc_hd__a221oi_1 _11279_ (.A1(net1073),
    .A2(_01322_),
    .B1(_01934_),
    .B2(net1249),
    .C1(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__a22oi_1 _11280_ (.A1(net1171),
    .A2(_02247_),
    .B1(_02400_),
    .B2(net251),
    .Y(_05304_));
 sky130_fd_sc_hd__a22oi_1 _11281_ (.A1(net505),
    .A2(_01553_),
    .B1(_02327_),
    .B2(net233),
    .Y(_05305_));
 sky130_fd_sc_hd__nand3_1 _11282_ (.A(_05303_),
    .B(_05304_),
    .C(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__o22a_2 _11283_ (.A1(net387),
    .A2(_01170_),
    .B1(_05301_),
    .B2(_05306_),
    .X(\w_CPU_dmem_rd_data_a4[1] ));
 sky130_fd_sc_hd__a21oi_1 _11284_ (.A1(\CPU_Dmem_value_a5[6][20] ),
    .A2(_02172_),
    .B1(net101),
    .Y(_05307_));
 sky130_fd_sc_hd__a22oi_1 _11285_ (.A1(\CPU_Dmem_value_a5[14][20] ),
    .A2(_01631_),
    .B1(_01705_),
    .B2(\CPU_Dmem_value_a5[15][20] ),
    .Y(_05308_));
 sky130_fd_sc_hd__a22oi_1 _11286_ (.A1(\CPU_Dmem_value_a5[1][20] ),
    .A2(net73),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][20] ),
    .Y(_05309_));
 sky130_fd_sc_hd__a22oi_1 _11287_ (.A1(\CPU_Dmem_value_a5[10][20] ),
    .A2(_01322_),
    .B1(_01553_),
    .B2(\CPU_Dmem_value_a5[13][20] ),
    .Y(_05310_));
 sky130_fd_sc_hd__nand4_1 _11288_ (.A(_05307_),
    .B(_05308_),
    .C(_05309_),
    .D(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__a22o_1 _11289_ (.A1(\CPU_Dmem_value_a5[4][20] ),
    .A2(net54),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][20] ),
    .X(_05312_));
 sky130_fd_sc_hd__a221oi_1 _11290_ (.A1(\CPU_Dmem_value_a5[2][20] ),
    .A2(net65),
    .B1(net63),
    .B2(\CPU_Dmem_value_a5[3][20] ),
    .C1(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__a22oi_1 _11291_ (.A1(\CPU_Dmem_value_a5[12][20] ),
    .A2(net80),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][20] ),
    .Y(_05314_));
 sky130_fd_sc_hd__a22oi_1 _11292_ (.A1(\CPU_Dmem_value_a5[11][20] ),
    .A2(_01397_),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][20] ),
    .Y(_05315_));
 sky130_fd_sc_hd__nand3_1 _11293_ (.A(_05313_),
    .B(_05314_),
    .C(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o22a_1 _11294_ (.A1(net646),
    .A2(_01170_),
    .B1(_05311_),
    .B2(_05316_),
    .X(\w_CPU_dmem_rd_data_a4[20] ));
 sky130_fd_sc_hd__a21oi_1 _11295_ (.A1(net636),
    .A2(_02247_),
    .B1(net100),
    .Y(_05317_));
 sky130_fd_sc_hd__a22oi_1 _11296_ (.A1(net680),
    .A2(_01397_),
    .B1(_01705_),
    .B2(net982),
    .Y(_05318_));
 sky130_fd_sc_hd__a22oi_1 _11297_ (.A1(net476),
    .A2(net80),
    .B1(_02172_),
    .B2(net208),
    .Y(_05319_));
 sky130_fd_sc_hd__a22oi_1 _11298_ (.A1(net876),
    .A2(_01553_),
    .B1(net65),
    .B2(net577),
    .Y(_05320_));
 sky130_fd_sc_hd__nand4_1 _11299_ (.A(_05317_),
    .B(_05318_),
    .C(_05319_),
    .D(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__a22oi_1 _11300_ (.A1(net575),
    .A2(_01631_),
    .B1(_02400_),
    .B2(net1042),
    .Y(_05322_));
 sky130_fd_sc_hd__a22oi_1 _11301_ (.A1(net277),
    .A2(net62),
    .B1(net43),
    .B2(net403),
    .Y(_05323_));
 sky130_fd_sc_hd__a22oi_1 _11302_ (.A1(net799),
    .A2(net72),
    .B1(net55),
    .B2(net686),
    .Y(_05324_));
 sky130_fd_sc_hd__a22oi_1 _11303_ (.A1(net349),
    .A2(_01322_),
    .B1(_02092_),
    .B2(net765),
    .Y(_05325_));
 sky130_fd_sc_hd__nand4_1 _11304_ (.A(_05322_),
    .B(_05323_),
    .C(_05324_),
    .D(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__o22a_1 _11305_ (.A1(net838),
    .A2(_01170_),
    .B1(_05321_),
    .B2(_05326_),
    .X(\w_CPU_dmem_rd_data_a4[21] ));
 sky130_fd_sc_hd__a21oi_1 _11306_ (.A1(net747),
    .A2(_02172_),
    .B1(net100),
    .Y(_05327_));
 sky130_fd_sc_hd__a22oi_1 _11307_ (.A1(\CPU_Dmem_value_a5[12][22] ),
    .A2(net81),
    .B1(_01631_),
    .B2(\CPU_Dmem_value_a5[14][22] ),
    .Y(_05328_));
 sky130_fd_sc_hd__a22oi_1 _11308_ (.A1(\CPU_Dmem_value_a5[13][22] ),
    .A2(_01553_),
    .B1(net55),
    .B2(\CPU_Dmem_value_a5[4][22] ),
    .Y(_05329_));
 sky130_fd_sc_hd__a22oi_1 _11309_ (.A1(\CPU_Dmem_value_a5[15][22] ),
    .A2(_01705_),
    .B1(net64),
    .B2(net1753),
    .Y(_05330_));
 sky130_fd_sc_hd__nand4_1 _11310_ (.A(_05327_),
    .B(_05328_),
    .C(_05329_),
    .D(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a22o_1 _11311_ (.A1(\CPU_Dmem_value_a5[5][22] ),
    .A2(_02092_),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][22] ),
    .X(_05332_));
 sky130_fd_sc_hd__a221oi_2 _11312_ (.A1(\CPU_Dmem_value_a5[1][22] ),
    .A2(net72),
    .B1(net62),
    .B2(\CPU_Dmem_value_a5[3][22] ),
    .C1(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__a22oi_1 _11313_ (.A1(\CPU_Dmem_value_a5[11][22] ),
    .A2(_01397_),
    .B1(net43),
    .B2(\CPU_Dmem_value_a5[8][22] ),
    .Y(_05334_));
 sky130_fd_sc_hd__a22oi_1 _11314_ (.A1(\CPU_Dmem_value_a5[10][22] ),
    .A2(_01322_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][22] ),
    .Y(_05335_));
 sky130_fd_sc_hd__nand3_1 _11315_ (.A(_05333_),
    .B(_05334_),
    .C(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__o22a_1 _11316_ (.A1(net1077),
    .A2(_01170_),
    .B1(net1754),
    .B2(_05336_),
    .X(\w_CPU_dmem_rd_data_a4[22] ));
 sky130_fd_sc_hd__a21oi_1 _11317_ (.A1(\CPU_Dmem_value_a5[4][23] ),
    .A2(net54),
    .B1(net101),
    .Y(_05337_));
 sky130_fd_sc_hd__a22oi_1 _11318_ (.A1(\CPU_Dmem_value_a5[10][23] ),
    .A2(_01322_),
    .B1(net65),
    .B2(\CPU_Dmem_value_a5[2][23] ),
    .Y(_05338_));
 sky130_fd_sc_hd__a22oi_1 _11319_ (.A1(\CPU_Dmem_value_a5[12][23] ),
    .A2(_01478_),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][23] ),
    .Y(_05339_));
 sky130_fd_sc_hd__a22oi_1 _11320_ (.A1(\CPU_Dmem_value_a5[14][23] ),
    .A2(_01631_),
    .B1(net73),
    .B2(\CPU_Dmem_value_a5[1][23] ),
    .Y(_05340_));
 sky130_fd_sc_hd__nand4_1 _11321_ (.A(_05337_),
    .B(_05338_),
    .C(_05339_),
    .D(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__a22o_1 _11322_ (.A1(\CPU_Dmem_value_a5[3][23] ),
    .A2(net63),
    .B1(net44),
    .B2(\CPU_Dmem_value_a5[8][23] ),
    .X(_05342_));
 sky130_fd_sc_hd__a221oi_1 _11323_ (.A1(\CPU_Dmem_value_a5[15][23] ),
    .A2(_01705_),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][23] ),
    .C1(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__a22oi_1 _11324_ (.A1(\CPU_Dmem_value_a5[13][23] ),
    .A2(_01553_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][23] ),
    .Y(_05344_));
 sky130_fd_sc_hd__a22oi_1 _11325_ (.A1(\CPU_Dmem_value_a5[11][23] ),
    .A2(_01397_),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][23] ),
    .Y(_05345_));
 sky130_fd_sc_hd__nand3_1 _11326_ (.A(_05343_),
    .B(_05344_),
    .C(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__o22a_1 _11327_ (.A1(net775),
    .A2(_01170_),
    .B1(_05341_),
    .B2(_05346_),
    .X(\w_CPU_dmem_rd_data_a4[23] ));
 sky130_fd_sc_hd__a21oi_1 _11328_ (.A1(net363),
    .A2(_02092_),
    .B1(net100),
    .Y(_05347_));
 sky130_fd_sc_hd__a22oi_1 _11329_ (.A1(net781),
    .A2(_01631_),
    .B1(net62),
    .B2(net231),
    .Y(_05348_));
 sky130_fd_sc_hd__a22oi_1 _11330_ (.A1(net468),
    .A2(net64),
    .B1(_02247_),
    .B2(net581),
    .Y(_05349_));
 sky130_fd_sc_hd__a22oi_1 _11331_ (.A1(\CPU_Dmem_value_a5[11][24] ),
    .A2(_01397_),
    .B1(_01705_),
    .B2(net293),
    .Y(_05350_));
 sky130_fd_sc_hd__nand4_1 _11332_ (.A(_05347_),
    .B(_05348_),
    .C(_05349_),
    .D(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a22o_1 _11333_ (.A1(\CPU_Dmem_value_a5[4][24] ),
    .A2(net54),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][24] ),
    .X(_05352_));
 sky130_fd_sc_hd__a221oi_1 _11334_ (.A1(\CPU_Dmem_value_a5[12][24] ),
    .A2(net81),
    .B1(net73),
    .B2(\CPU_Dmem_value_a5[1][24] ),
    .C1(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__a22oi_1 _11335_ (.A1(\CPU_Dmem_value_a5[10][24] ),
    .A2(_01322_),
    .B1(_02400_),
    .B2(net1708),
    .Y(_05354_));
 sky130_fd_sc_hd__a22oi_1 _11336_ (.A1(\CPU_Dmem_value_a5[13][24] ),
    .A2(_01553_),
    .B1(net43),
    .B2(\CPU_Dmem_value_a5[8][24] ),
    .Y(_05355_));
 sky130_fd_sc_hd__nand3_1 _11337_ (.A(_05353_),
    .B(_05354_),
    .C(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__o22a_2 _11338_ (.A1(net383),
    .A2(_01170_),
    .B1(_05351_),
    .B2(_05356_),
    .X(\w_CPU_dmem_rd_data_a4[24] ));
 sky130_fd_sc_hd__a21oi_1 _11339_ (.A1(net265),
    .A2(net44),
    .B1(net100),
    .Y(_05357_));
 sky130_fd_sc_hd__a22oi_1 _11340_ (.A1(\CPU_Dmem_value_a5[10][25] ),
    .A2(_01322_),
    .B1(_02092_),
    .B2(net797),
    .Y(_05358_));
 sky130_fd_sc_hd__a22oi_1 _11341_ (.A1(\CPU_Dmem_value_a5[1][25] ),
    .A2(net72),
    .B1(_02247_),
    .B2(net440),
    .Y(_05359_));
 sky130_fd_sc_hd__a22oi_1 _11342_ (.A1(net1057),
    .A2(_01397_),
    .B1(net81),
    .B2(net253),
    .Y(_05360_));
 sky130_fd_sc_hd__nand4_1 _11343_ (.A(_05357_),
    .B(_05358_),
    .C(_05359_),
    .D(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__a22o_1 _11344_ (.A1(\CPU_Dmem_value_a5[4][25] ),
    .A2(net54),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][25] ),
    .X(_05362_));
 sky130_fd_sc_hd__a221oi_1 _11345_ (.A1(net1012),
    .A2(_01631_),
    .B1(net63),
    .B2(net1020),
    .C1(_05362_),
    .Y(_05363_));
 sky130_fd_sc_hd__a22oi_1 _11346_ (.A1(\CPU_Dmem_value_a5[15][25] ),
    .A2(_01705_),
    .B1(net64),
    .B2(net301),
    .Y(_05364_));
 sky130_fd_sc_hd__a22oi_1 _11347_ (.A1(net365),
    .A2(_01553_),
    .B1(_02400_),
    .B2(net545),
    .Y(_05365_));
 sky130_fd_sc_hd__nand3_1 _11348_ (.A(_05363_),
    .B(_05364_),
    .C(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__o22a_2 _11349_ (.A1(net553),
    .A2(_01170_),
    .B1(_05361_),
    .B2(_05366_),
    .X(\w_CPU_dmem_rd_data_a4[25] ));
 sky130_fd_sc_hd__a21oi_1 _11350_ (.A1(net610),
    .A2(net72),
    .B1(net99),
    .Y(_05367_));
 sky130_fd_sc_hd__a22oi_1 _11351_ (.A1(\CPU_Dmem_value_a5[10][26] ),
    .A2(_01322_),
    .B1(_01553_),
    .B2(\CPU_Dmem_value_a5[13][26] ),
    .Y(_05368_));
 sky130_fd_sc_hd__a22oi_1 _11352_ (.A1(\CPU_Dmem_value_a5[15][26] ),
    .A2(_01705_),
    .B1(net62),
    .B2(\CPU_Dmem_value_a5[3][26] ),
    .Y(_05369_));
 sky130_fd_sc_hd__a22oi_1 _11353_ (.A1(\CPU_Dmem_value_a5[11][26] ),
    .A2(_01397_),
    .B1(net64),
    .B2(\CPU_Dmem_value_a5[2][26] ),
    .Y(_05370_));
 sky130_fd_sc_hd__nand4_1 _11354_ (.A(_05367_),
    .B(_05368_),
    .C(_05369_),
    .D(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__a22oi_1 _11355_ (.A1(net511),
    .A2(_02247_),
    .B1(_02400_),
    .B2(net429),
    .Y(_05372_));
 sky130_fd_sc_hd__a22oi_1 _11356_ (.A1(net281),
    .A2(net55),
    .B1(net43),
    .B2(net972),
    .Y(_05373_));
 sky130_fd_sc_hd__a22oi_1 _11357_ (.A1(net880),
    .A2(net81),
    .B1(_01631_),
    .B2(net257),
    .Y(_05374_));
 sky130_fd_sc_hd__a22oi_1 _11358_ (.A1(net915),
    .A2(_02092_),
    .B1(_02172_),
    .B2(net668),
    .Y(_05375_));
 sky130_fd_sc_hd__nand4_1 _11359_ (.A(_05372_),
    .B(_05373_),
    .C(_05374_),
    .D(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__o22a_1 _11360_ (.A1(net1075),
    .A2(_01170_),
    .B1(_05371_),
    .B2(_05376_),
    .X(\w_CPU_dmem_rd_data_a4[26] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__a21oi_1 _11362_ (.A1(net852),
    .A2(net43),
    .B1(net99),
    .Y(_05378_));
 sky130_fd_sc_hd__a22oi_1 _11363_ (.A1(net850),
    .A2(_01322_),
    .B1(_02247_),
    .B2(net215),
    .Y(_05379_));
 sky130_fd_sc_hd__a22oi_1 _11364_ (.A1(net896),
    .A2(_01397_),
    .B1(net62),
    .B2(net1067),
    .Y(_05380_));
 sky130_fd_sc_hd__a22oi_1 _11365_ (.A1(net589),
    .A2(_01631_),
    .B1(net64),
    .B2(net397),
    .Y(_05381_));
 sky130_fd_sc_hd__nand4_1 _11366_ (.A(_05378_),
    .B(_05379_),
    .C(_05380_),
    .D(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__a22o_1 _11367_ (.A1(net1254),
    .A2(net55),
    .B1(_02092_),
    .B2(net1273),
    .X(_05383_));
 sky130_fd_sc_hd__a221oi_1 _11368_ (.A1(net815),
    .A2(_01553_),
    .B1(_02172_),
    .B2(net862),
    .C1(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__a22oi_1 _11369_ (.A1(net452),
    .A2(net81),
    .B1(net72),
    .B2(net389),
    .Y(_05385_));
 sky130_fd_sc_hd__a22oi_1 _11370_ (.A1(net425),
    .A2(_01705_),
    .B1(_02400_),
    .B2(net836),
    .Y(_05386_));
 sky130_fd_sc_hd__nand3_1 _11371_ (.A(_05384_),
    .B(_05385_),
    .C(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__o22a_1 _11372_ (.A1(net844),
    .A2(_01170_),
    .B1(_05382_),
    .B2(_05387_),
    .X(\w_CPU_dmem_rd_data_a4[27] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__a21oi_1 _11374_ (.A1(net648),
    .A2(_02247_),
    .B1(net99),
    .Y(_05389_));
 sky130_fd_sc_hd__a22oi_1 _11375_ (.A1(net1014),
    .A2(_01553_),
    .B1(_02172_),
    .B2(net415),
    .Y(_05390_));
 sky130_fd_sc_hd__a22oi_1 _11376_ (.A1(net442),
    .A2(_01397_),
    .B1(net64),
    .B2(net703),
    .Y(_05391_));
 sky130_fd_sc_hd__a22oi_1 _11377_ (.A1(net984),
    .A2(_01322_),
    .B1(_01705_),
    .B2(net217),
    .Y(_05392_));
 sky130_fd_sc_hd__nand4_1 _11378_ (.A(_05389_),
    .B(_05390_),
    .C(_05391_),
    .D(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__a22o_1 _11379_ (.A1(\CPU_Dmem_value_a5[4][28] ),
    .A2(net55),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][28] ),
    .X(_05394_));
 sky130_fd_sc_hd__a221oi_1 _11380_ (.A1(net938),
    .A2(net72),
    .B1(net62),
    .B2(net444),
    .C1(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__a22oi_1 _11381_ (.A1(net713),
    .A2(_01631_),
    .B1(net43),
    .B2(net886),
    .Y(_05396_));
 sky130_fd_sc_hd__a22oi_1 _11382_ (.A1(net823),
    .A2(net81),
    .B1(_02400_),
    .B2(net795),
    .Y(_05397_));
 sky130_fd_sc_hd__nand3_1 _11383_ (.A(_05395_),
    .B(_05396_),
    .C(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o22a_1 _11384_ (.A1(net753),
    .A2(_01170_),
    .B1(_05393_),
    .B2(_05398_),
    .X(\w_CPU_dmem_rd_data_a4[28] ));
 sky130_fd_sc_hd__a21oi_1 _11385_ (.A1(net259),
    .A2(net44),
    .B1(net100),
    .Y(_05399_));
 sky130_fd_sc_hd__a22oi_1 _11386_ (.A1(\CPU_Dmem_value_a5[11][29] ),
    .A2(_01397_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][29] ),
    .Y(_05400_));
 sky130_fd_sc_hd__a22oi_1 _11387_ (.A1(\CPU_Dmem_value_a5[12][29] ),
    .A2(net80),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][29] ),
    .Y(_05401_));
 sky130_fd_sc_hd__a22oi_1 _11388_ (.A1(\CPU_Dmem_value_a5[14][29] ),
    .A2(_01631_),
    .B1(net72),
    .B2(\CPU_Dmem_value_a5[1][29] ),
    .Y(_05402_));
 sky130_fd_sc_hd__nand4_1 _11389_ (.A(_05399_),
    .B(_05400_),
    .C(_05401_),
    .D(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a22o_1 _11390_ (.A1(\CPU_Dmem_value_a5[4][29] ),
    .A2(net54),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][29] ),
    .X(_05404_));
 sky130_fd_sc_hd__a221oi_1 _11391_ (.A1(\CPU_Dmem_value_a5[13][29] ),
    .A2(_01553_),
    .B1(net63),
    .B2(net1821),
    .C1(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__a22oi_1 _11392_ (.A1(\CPU_Dmem_value_a5[10][29] ),
    .A2(_01322_),
    .B1(_01705_),
    .B2(\CPU_Dmem_value_a5[15][29] ),
    .Y(_05406_));
 sky130_fd_sc_hd__a22oi_1 _11393_ (.A1(\CPU_Dmem_value_a5[2][29] ),
    .A2(net65),
    .B1(_02172_),
    .B2(\CPU_Dmem_value_a5[6][29] ),
    .Y(_05407_));
 sky130_fd_sc_hd__nand3_1 _11394_ (.A(_05405_),
    .B(_05406_),
    .C(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__o22a_1 _11395_ (.A1(net369),
    .A2(_01170_),
    .B1(_05403_),
    .B2(_05408_),
    .X(\w_CPU_dmem_rd_data_a4[29] ));
 sky130_fd_sc_hd__a21oi_1 _11396_ (.A1(net1071),
    .A2(_02018_),
    .B1(_01177_),
    .Y(_05409_));
 sky130_fd_sc_hd__a22oi_1 _11397_ (.A1(net466),
    .A2(_01322_),
    .B1(_01934_),
    .B2(net1107),
    .Y(_05410_));
 sky130_fd_sc_hd__a22oi_1 _11398_ (.A1(net1348),
    .A2(_01553_),
    .B1(_02172_),
    .B2(net1032),
    .Y(_05411_));
 sky130_fd_sc_hd__a22oi_1 _11399_ (.A1(net1219),
    .A2(_01478_),
    .B1(_01782_),
    .B2(net690),
    .Y(_05412_));
 sky130_fd_sc_hd__nand4_1 _11400_ (.A(_05409_),
    .B(_05410_),
    .C(_05411_),
    .D(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__a22o_1 _11401_ (.A1(net1004),
    .A2(_01861_),
    .B1(_02400_),
    .B2(net1341),
    .X(_05414_));
 sky130_fd_sc_hd__a221oi_1 _11402_ (.A1(net805),
    .A2(_01397_),
    .B1(_01705_),
    .B2(net1316),
    .C1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__a22oi_1 _11403_ (.A1(net1191),
    .A2(_02092_),
    .B1(_02247_),
    .B2(net1079),
    .Y(_05416_));
 sky130_fd_sc_hd__a22oi_1 _11404_ (.A1(net1221),
    .A2(_01631_),
    .B1(_02327_),
    .B2(net626),
    .Y(_05417_));
 sky130_fd_sc_hd__nand3_1 _11405_ (.A(_05415_),
    .B(_05416_),
    .C(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__o22a_1 _11406_ (.A1(net399),
    .A2(_01170_),
    .B1(_05413_),
    .B2(_05418_),
    .X(\w_CPU_dmem_rd_data_a4[2] ));
 sky130_fd_sc_hd__a21oi_1 _11407_ (.A1(net263),
    .A2(net55),
    .B1(net99),
    .Y(_05419_));
 sky130_fd_sc_hd__a22oi_1 _11408_ (.A1(net682),
    .A2(net81),
    .B1(_01553_),
    .B2(net1046),
    .Y(_05420_));
 sky130_fd_sc_hd__a22oi_1 _11409_ (.A1(net482),
    .A2(_01322_),
    .B1(_02172_),
    .B2(net727),
    .Y(_05421_));
 sky130_fd_sc_hd__a22oi_1 _11410_ (.A1(net407),
    .A2(_01397_),
    .B1(_01631_),
    .B2(net996),
    .Y(_05422_));
 sky130_fd_sc_hd__nand4_1 _11411_ (.A(_05419_),
    .B(_05420_),
    .C(_05421_),
    .D(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__a22o_1 _11412_ (.A1(net773),
    .A2(net64),
    .B1(_02400_),
    .B2(net210),
    .X(_05424_));
 sky130_fd_sc_hd__a221oi_1 _11413_ (.A1(net858),
    .A2(_01705_),
    .B1(net62),
    .B2(net944),
    .C1(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__a22oi_1 _11414_ (.A1(net769),
    .A2(_02092_),
    .B1(_02247_),
    .B2(net1090),
    .Y(_05426_));
 sky130_fd_sc_hd__a22oi_1 _11415_ (.A1(net644),
    .A2(net72),
    .B1(net43),
    .B2(net892),
    .Y(_05427_));
 sky130_fd_sc_hd__nand3_1 _11416_ (.A(_05425_),
    .B(_05426_),
    .C(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__o22a_1 _11417_ (.A1(net1083),
    .A2(_01170_),
    .B1(_05423_),
    .B2(_05428_),
    .X(\w_CPU_dmem_rd_data_a4[30] ));
 sky130_fd_sc_hd__a22oi_1 _11418_ (.A1(net903),
    .A2(_01322_),
    .B1(_02400_),
    .B2(net634),
    .Y(_05429_));
 sky130_fd_sc_hd__a22oi_1 _11419_ (.A1(net1132),
    .A2(_01705_),
    .B1(net72),
    .B2(net297),
    .Y(_05430_));
 sky130_fd_sc_hd__a22oi_1 _11420_ (.A1(net913),
    .A2(_01553_),
    .B1(net65),
    .B2(net1026),
    .Y(_05431_));
 sky130_fd_sc_hd__a22oi_1 _11421_ (.A1(net1116),
    .A2(net62),
    .B1(_02092_),
    .B2(net1006),
    .Y(_05432_));
 sky130_fd_sc_hd__nand4_1 _11422_ (.A(_05429_),
    .B(_05430_),
    .C(_05431_),
    .D(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__mux2i_1 _11423_ (.A0(\CPU_Dmem_value_a5[4][31] ),
    .A1(\CPU_Dmem_value_a5[12][31] ),
    .S(\CPU_dmem_addr_a4[3] ),
    .Y(_05434_));
 sky130_fd_sc_hd__o21ai_0 _11424_ (.A1(\CPU_Dmem_value_a5[8][31] ),
    .A2(_01317_),
    .B1(_01166_),
    .Y(_05435_));
 sky130_fd_sc_hd__a21oi_2 _11425_ (.A1(\CPU_dmem_addr_a4[2] ),
    .A2(_05434_),
    .B1(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__a22oi_1 _11426_ (.A1(net1044),
    .A2(_01631_),
    .B1(_02247_),
    .B2(net283),
    .Y(_05437_));
 sky130_fd_sc_hd__a22oi_1 _11427_ (.A1(net620),
    .A2(_01397_),
    .B1(_02172_),
    .B2(net287),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _11428_ (.A(_05437_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__o32a_1 _11429_ (.A1(_05433_),
    .A2(_05436_),
    .A3(_05439_),
    .B1(_01170_),
    .B2(net450),
    .X(\w_CPU_dmem_rd_data_a4[31] ));
 sky130_fd_sc_hd__a21oi_1 _11430_ (.A1(net513),
    .A2(_01861_),
    .B1(_01177_),
    .Y(_05440_));
 sky130_fd_sc_hd__a22oi_1 _11431_ (.A1(net1231),
    .A2(_01478_),
    .B1(_01782_),
    .B2(net565),
    .Y(_05441_));
 sky130_fd_sc_hd__a22oi_1 _11432_ (.A1(net642),
    .A2(_02172_),
    .B1(_02400_),
    .B2(net1321),
    .Y(_05442_));
 sky130_fd_sc_hd__a22oi_1 _11433_ (.A1(net1127),
    .A2(_01322_),
    .B1(_01397_),
    .B2(net1059),
    .Y(_05443_));
 sky130_fd_sc_hd__nand4_1 _11434_ (.A(_05440_),
    .B(_05441_),
    .C(_05442_),
    .D(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__a22o_1 _11435_ (.A1(\CPU_Dmem_value_a5[3][3] ),
    .A2(_01934_),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][3] ),
    .X(_05445_));
 sky130_fd_sc_hd__a221oi_1 _11436_ (.A1(net1264),
    .A2(_01553_),
    .B1(_02018_),
    .B2(net830),
    .C1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__a22oi_1 _11437_ (.A1(net1053),
    .A2(_01705_),
    .B1(_02247_),
    .B2(net749),
    .Y(_05447_));
 sky130_fd_sc_hd__a22oi_1 _11438_ (.A1(net1257),
    .A2(_01631_),
    .B1(_02327_),
    .B2(net1160),
    .Y(_05448_));
 sky130_fd_sc_hd__nand3_1 _11439_ (.A(_05446_),
    .B(_05447_),
    .C(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__o22a_1 _11440_ (.A1(net992),
    .A2(_01170_),
    .B1(_05444_),
    .B2(_05449_),
    .X(\w_CPU_dmem_rd_data_a4[3] ));
 sky130_fd_sc_hd__a21oi_1 _11441_ (.A1(net419),
    .A2(_02400_),
    .B1(net101),
    .Y(_05450_));
 sky130_fd_sc_hd__a22oi_1 _11442_ (.A1(net745),
    .A2(_01397_),
    .B1(_01631_),
    .B2(net212),
    .Y(_05451_));
 sky130_fd_sc_hd__a22oi_1 _11443_ (.A1(\CPU_Dmem_value_a5[1][4] ),
    .A2(_01782_),
    .B1(_02172_),
    .B2(net235),
    .Y(_05452_));
 sky130_fd_sc_hd__a22oi_1 _11444_ (.A1(net920),
    .A2(_01322_),
    .B1(_01478_),
    .B2(net517),
    .Y(_05453_));
 sky130_fd_sc_hd__nand4_1 _11445_ (.A(_05450_),
    .B(_05451_),
    .C(_05452_),
    .D(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a22o_1 _11446_ (.A1(\CPU_Dmem_value_a5[4][4] ),
    .A2(_02018_),
    .B1(_02092_),
    .B2(\CPU_Dmem_value_a5[5][4] ),
    .X(_05455_));
 sky130_fd_sc_hd__a221oi_1 _11447_ (.A1(net484),
    .A2(_01861_),
    .B1(net63),
    .B2(net327),
    .C1(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__a22oi_1 _11448_ (.A1(net654),
    .A2(_01553_),
    .B1(net44),
    .B2(net337),
    .Y(_05457_));
 sky130_fd_sc_hd__a22oi_1 _11449_ (.A1(net509),
    .A2(_01705_),
    .B1(_02247_),
    .B2(net502),
    .Y(_05458_));
 sky130_fd_sc_hd__nand3_1 _11450_ (.A(_05456_),
    .B(_05457_),
    .C(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__o22a_2 _11451_ (.A1(net729),
    .A2(_01170_),
    .B1(_05454_),
    .B2(_05459_),
    .X(\w_CPU_dmem_rd_data_a4[4] ));
 sky130_fd_sc_hd__a21oi_1 _11452_ (.A1(net832),
    .A2(_02400_),
    .B1(_01177_),
    .Y(_05460_));
 sky130_fd_sc_hd__a22oi_1 _11453_ (.A1(net1344),
    .A2(_01478_),
    .B1(_01861_),
    .B2(net1199),
    .Y(_05461_));
 sky130_fd_sc_hd__a22oi_1 _11454_ (.A1(net860),
    .A2(_01934_),
    .B1(_02092_),
    .B2(net1097),
    .Y(_05462_));
 sky130_fd_sc_hd__a22oi_1 _11455_ (.A1(net361),
    .A2(_01322_),
    .B1(_01631_),
    .B2(net427),
    .Y(_05463_));
 sky130_fd_sc_hd__nand4_1 _11456_ (.A(_05460_),
    .B(_05461_),
    .C(_05462_),
    .D(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__a22oi_1 _11457_ (.A1(net1174),
    .A2(_01397_),
    .B1(_02018_),
    .B2(net1040),
    .Y(_05465_));
 sky130_fd_sc_hd__a22oi_1 _11458_ (.A1(net954),
    .A2(_01705_),
    .B1(_02327_),
    .B2(net1166),
    .Y(_05466_));
 sky130_fd_sc_hd__a22oi_1 _11459_ (.A1(net958),
    .A2(_01782_),
    .B1(_02172_),
    .B2(net956),
    .Y(_05467_));
 sky130_fd_sc_hd__a22oi_1 _11460_ (.A1(net994),
    .A2(_01553_),
    .B1(_02247_),
    .B2(net591),
    .Y(_05468_));
 sky130_fd_sc_hd__nand4_1 _11461_ (.A(_05465_),
    .B(_05466_),
    .C(_05467_),
    .D(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__o22a_1 _11462_ (.A1(net488),
    .A2(_01170_),
    .B1(_05464_),
    .B2(_05469_),
    .X(\w_CPU_dmem_rd_data_a4[5] ));
 sky130_fd_sc_hd__a21oi_1 _11463_ (.A1(net1123),
    .A2(_02247_),
    .B1(net99),
    .Y(_05470_));
 sky130_fd_sc_hd__a22oi_1 _11464_ (.A1(net1202),
    .A2(net81),
    .B1(_01553_),
    .B2(net291),
    .Y(_05471_));
 sky130_fd_sc_hd__a22oi_1 _11465_ (.A1(net705),
    .A2(_01631_),
    .B1(net72),
    .B2(net976),
    .Y(_05472_));
 sky130_fd_sc_hd__a22oi_1 _11466_ (.A1(net950),
    .A2(_01322_),
    .B1(net55),
    .B2(net1158),
    .Y(_05473_));
 sky130_fd_sc_hd__nand4_1 _11467_ (.A(_05470_),
    .B(_05471_),
    .C(_05472_),
    .D(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(\CPU_Dmem_value_a5[3][6] ),
    .A2(net62),
    .B1(_02092_),
    .B2(net1422),
    .X(_05475_));
 sky130_fd_sc_hd__a221oi_1 _11469_ (.A1(net755),
    .A2(net64),
    .B1(_02172_),
    .B2(net907),
    .C1(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__a22oi_1 _11470_ (.A1(net630),
    .A2(_01397_),
    .B1(net43),
    .B2(net811),
    .Y(_05477_));
 sky130_fd_sc_hd__a22oi_1 _11471_ (.A1(net1143),
    .A2(_01705_),
    .B1(_02400_),
    .B2(net898),
    .Y(_05478_));
 sky130_fd_sc_hd__nand3_1 _11472_ (.A(_05476_),
    .B(_05477_),
    .C(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__o22a_1 _11473_ (.A1(net890),
    .A2(_01170_),
    .B1(_05474_),
    .B2(_05479_),
    .X(\w_CPU_dmem_rd_data_a4[6] ));
 sky130_fd_sc_hd__a21oi_1 _11474_ (.A1(net587),
    .A2(net44),
    .B1(net101),
    .Y(_05480_));
 sky130_fd_sc_hd__a22oi_1 _11475_ (.A1(\CPU_Dmem_value_a5[15][7] ),
    .A2(_01705_),
    .B1(_02400_),
    .B2(\CPU_Dmem_value_a5[9][7] ),
    .Y(_05481_));
 sky130_fd_sc_hd__a22oi_1 _11476_ (.A1(\CPU_Dmem_value_a5[10][7] ),
    .A2(_01322_),
    .B1(net65),
    .B2(net854),
    .Y(_05482_));
 sky130_fd_sc_hd__a22oi_1 _11477_ (.A1(net968),
    .A2(_01397_),
    .B1(_01553_),
    .B2(net678),
    .Y(_05483_));
 sky130_fd_sc_hd__nand4_1 _11478_ (.A(_05480_),
    .B(_05481_),
    .C(_05482_),
    .D(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__a22o_1 _11479_ (.A1(\CPU_Dmem_value_a5[3][7] ),
    .A2(net63),
    .B1(net54),
    .B2(\CPU_Dmem_value_a5[4][7] ),
    .X(_05485_));
 sky130_fd_sc_hd__a221oi_1 _11480_ (.A1(net868),
    .A2(_01782_),
    .B1(_02172_),
    .B2(net507),
    .C1(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__a22oi_1 _11481_ (.A1(\CPU_Dmem_value_a5[12][7] ),
    .A2(_01478_),
    .B1(_02092_),
    .B2(net652),
    .Y(_05487_));
 sky130_fd_sc_hd__a22oi_1 _11482_ (.A1(net319),
    .A2(_01631_),
    .B1(_02247_),
    .B2(net317),
    .Y(_05488_));
 sky130_fd_sc_hd__nand3_1 _11483_ (.A(_05486_),
    .B(_05487_),
    .C(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__o22a_1 _11484_ (.A1(net789),
    .A2(_01170_),
    .B1(_05484_),
    .B2(_05489_),
    .X(\w_CPU_dmem_rd_data_a4[7] ));
 sky130_fd_sc_hd__a21oi_1 _11485_ (.A1(net771),
    .A2(_02092_),
    .B1(_01177_),
    .Y(_05490_));
 sky130_fd_sc_hd__a22oi_1 _11486_ (.A1(net672),
    .A2(_01397_),
    .B1(_01782_),
    .B2(net525),
    .Y(_05491_));
 sky130_fd_sc_hd__a22oi_1 _11487_ (.A1(net725),
    .A2(_01705_),
    .B1(_01861_),
    .B2(net279),
    .Y(_05492_));
 sky130_fd_sc_hd__a22oi_1 _11488_ (.A1(net1700),
    .A2(_01553_),
    .B1(_01631_),
    .B2(net932),
    .Y(_05493_));
 sky130_fd_sc_hd__nand4_1 _11489_ (.A(_05490_),
    .B(_05491_),
    .C(_05492_),
    .D(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__a22o_1 _11490_ (.A1(\CPU_Dmem_value_a5[4][8] ),
    .A2(_02018_),
    .B1(_02247_),
    .B2(\CPU_Dmem_value_a5[7][8] ),
    .X(_05495_));
 sky130_fd_sc_hd__a221oi_1 _11491_ (.A1(net870),
    .A2(_01934_),
    .B1(_02172_),
    .B2(net842),
    .C1(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__a22oi_1 _11492_ (.A1(net492),
    .A2(_01322_),
    .B1(_02327_),
    .B2(net763),
    .Y(_05497_));
 sky130_fd_sc_hd__a22oi_1 _11493_ (.A1(net761),
    .A2(_01478_),
    .B1(_02400_),
    .B2(net658),
    .Y(_05498_));
 sky130_fd_sc_hd__nand3_1 _11494_ (.A(_05496_),
    .B(_05497_),
    .C(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__o22a_2 _11495_ (.A1(net539),
    .A2(_01170_),
    .B1(_05494_),
    .B2(_05499_),
    .X(\w_CPU_dmem_rd_data_a4[8] ));
 sky130_fd_sc_hd__a22oi_1 _11496_ (.A1(net1246),
    .A2(_01553_),
    .B1(_01631_),
    .B2(net988),
    .Y(_05500_));
 sky130_fd_sc_hd__a21oi_1 _11497_ (.A1(net1229),
    .A2(_02092_),
    .B1(net101),
    .Y(_05501_));
 sky130_fd_sc_hd__a22oi_1 _11498_ (.A1(net1697),
    .A2(net80),
    .B1(net63),
    .B2(net313),
    .Y(_05502_));
 sky130_fd_sc_hd__a22oi_1 _11499_ (.A1(\CPU_Dmem_value_a5[15][9] ),
    .A2(_01705_),
    .B1(_01782_),
    .B2(net707),
    .Y(_05503_));
 sky130_fd_sc_hd__nand4_1 _11500_ (.A(_05500_),
    .B(_05501_),
    .C(_05502_),
    .D(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__a22oi_1 _11501_ (.A1(net454),
    .A2(_01322_),
    .B1(_02400_),
    .B2(net1352),
    .Y(_05505_));
 sky130_fd_sc_hd__a22oi_1 _11502_ (.A1(net1362),
    .A2(_02018_),
    .B1(_02172_),
    .B2(net1630),
    .Y(_05506_));
 sky130_fd_sc_hd__a22oi_1 _11503_ (.A1(net1154),
    .A2(net65),
    .B1(net44),
    .B2(net470),
    .Y(_05507_));
 sky130_fd_sc_hd__a22oi_1 _11504_ (.A1(net1329),
    .A2(_01397_),
    .B1(_02247_),
    .B2(net379),
    .Y(_05508_));
 sky130_fd_sc_hd__nand4_1 _11505_ (.A(_05505_),
    .B(_05506_),
    .C(_05507_),
    .D(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__o22a_1 _11506_ (.A1(net1381),
    .A2(_01170_),
    .B1(net1698),
    .B2(_05509_),
    .X(\w_CPU_dmem_rd_data_a4[9] ));
 sky130_fd_sc_hd__fa_1 _11507_ (.A(_05510_),
    .B(_05511_),
    .CIN(_05512_),
    .COUT(_05513_),
    .SUM(_05514_));
 sky130_fd_sc_hd__fa_1 _11508_ (.A(_05511_),
    .B(_05515_),
    .CIN(_05516_),
    .COUT(_05517_),
    .SUM(_05518_));
 sky130_fd_sc_hd__fa_1 _11509_ (.A(_05519_),
    .B(_05520_),
    .CIN(_05521_),
    .COUT(_05522_),
    .SUM(\CPU_br_tgt_pc_a2[1] ));
 sky130_fd_sc_hd__ha_4 _11510_ (.A(_05523_),
    .B(\CPU_src2_value_a3[31] ),
    .COUT(_05524_),
    .SUM(_05525_));
 sky130_fd_sc_hd__ha_4 _11511_ (.A(_05526_),
    .B(\CPU_src2_value_a3[27] ),
    .COUT(_05527_),
    .SUM(_05528_));
 sky130_fd_sc_hd__ha_1 _11512_ (.A(\CPU_src1_value_a3[27] ),
    .B(\CPU_src2_value_a3[27] ),
    .COUT(_05529_),
    .SUM(_05530_));
 sky130_fd_sc_hd__ha_4 _11513_ (.A(_05531_),
    .B(\CPU_src2_value_a3[23] ),
    .COUT(_05532_),
    .SUM(_05533_));
 sky130_fd_sc_hd__ha_1 _11514_ (.A(\CPU_src1_value_a3[23] ),
    .B(\CPU_src2_value_a3[23] ),
    .COUT(_05534_),
    .SUM(_05535_));
 sky130_fd_sc_hd__ha_2 _11515_ (.A(_05536_),
    .B(\CPU_src2_value_a3[19] ),
    .COUT(_05537_),
    .SUM(_05538_));
 sky130_fd_sc_hd__ha_1 _11516_ (.A(\CPU_src1_value_a3[19] ),
    .B(\CPU_src2_value_a3[19] ),
    .COUT(_05539_),
    .SUM(_05540_));
 sky130_fd_sc_hd__ha_2 _11517_ (.A(_05541_),
    .B(\CPU_src2_value_a3[15] ),
    .COUT(_05542_),
    .SUM(_05543_));
 sky130_fd_sc_hd__ha_1 _11518_ (.A(\CPU_src1_value_a3[15] ),
    .B(\CPU_src2_value_a3[15] ),
    .COUT(_05544_),
    .SUM(_05545_));
 sky130_fd_sc_hd__ha_2 _11519_ (.A(_05546_),
    .B(\CPU_src2_value_a3[11] ),
    .COUT(_05547_),
    .SUM(_05548_));
 sky130_fd_sc_hd__ha_1 _11520_ (.A(\CPU_src1_value_a3[11] ),
    .B(\CPU_src2_value_a3[11] ),
    .COUT(_05549_),
    .SUM(_05550_));
 sky130_fd_sc_hd__ha_2 _11521_ (.A(_05551_),
    .B(\CPU_src2_value_a3[7] ),
    .COUT(_05552_),
    .SUM(_05553_));
 sky130_fd_sc_hd__ha_1 _11522_ (.A(\CPU_src1_value_a3[7] ),
    .B(\CPU_src2_value_a3[7] ),
    .COUT(_05554_),
    .SUM(_05555_));
 sky130_fd_sc_hd__ha_2 _11523_ (.A(_05556_),
    .B(\CPU_src2_value_a3[3] ),
    .COUT(_05557_),
    .SUM(_05558_));
 sky130_fd_sc_hd__ha_1 _11524_ (.A(\CPU_src1_value_a3[3] ),
    .B(\CPU_src2_value_a3[3] ),
    .COUT(_05559_),
    .SUM(_05560_));
 sky130_fd_sc_hd__ha_1 _11525_ (.A(_05511_),
    .B(\CPU_src2_value_a3[1] ),
    .COUT(_05561_),
    .SUM(_05562_));
 sky130_fd_sc_hd__ha_1 _11526_ (.A(\CPU_src1_value_a3[1] ),
    .B(\CPU_src2_value_a3[1] ),
    .COUT(_05563_),
    .SUM(_05564_));
 sky130_fd_sc_hd__ha_2 _11527_ (.A(\CPU_imm_a3[10] ),
    .B(_05565_),
    .COUT(_05566_),
    .SUM(_05567_));
 sky130_fd_sc_hd__ha_1 _11528_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[29] ),
    .COUT(_05568_),
    .SUM(_05569_));
 sky130_fd_sc_hd__ha_2 _11529_ (.A(\CPU_imm_a3[10] ),
    .B(_05570_),
    .COUT(_05571_),
    .SUM(_05572_));
 sky130_fd_sc_hd__ha_1 _11530_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[28] ),
    .COUT(_05573_),
    .SUM(_05574_));
 sky130_fd_sc_hd__ha_2 _11531_ (.A(\CPU_imm_a3[10] ),
    .B(_05526_),
    .COUT(_05575_),
    .SUM(_05576_));
 sky130_fd_sc_hd__ha_1 _11532_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[27] ),
    .COUT(_05577_),
    .SUM(_05578_));
 sky130_fd_sc_hd__ha_2 _11533_ (.A(\CPU_imm_a3[10] ),
    .B(_05579_),
    .COUT(_05580_),
    .SUM(_05581_));
 sky130_fd_sc_hd__ha_2 _11534_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[25] ),
    .COUT(_05582_),
    .SUM(_05583_));
 sky130_fd_sc_hd__ha_2 _11535_ (.A(\CPU_imm_a3[10] ),
    .B(_05584_),
    .COUT(_05585_),
    .SUM(_05586_));
 sky130_fd_sc_hd__ha_1 _11536_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[24] ),
    .COUT(_05587_),
    .SUM(_05588_));
 sky130_fd_sc_hd__ha_2 _11537_ (.A(\CPU_imm_a3[10] ),
    .B(_05531_),
    .COUT(_05589_),
    .SUM(_05590_));
 sky130_fd_sc_hd__ha_1 _11538_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[23] ),
    .COUT(_05591_),
    .SUM(_05592_));
 sky130_fd_sc_hd__ha_2 _11539_ (.A(\CPU_imm_a3[10] ),
    .B(_05536_),
    .COUT(_05593_),
    .SUM(_05594_));
 sky130_fd_sc_hd__ha_1 _11540_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[19] ),
    .COUT(_05595_),
    .SUM(_05596_));
 sky130_fd_sc_hd__ha_2 _11541_ (.A(\CPU_imm_a3[10] ),
    .B(_05597_),
    .COUT(_05598_),
    .SUM(_05599_));
 sky130_fd_sc_hd__ha_1 _11542_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[17] ),
    .COUT(_05600_),
    .SUM(_05601_));
 sky130_fd_sc_hd__ha_2 _11543_ (.A(\CPU_imm_a3[10] ),
    .B(_05602_),
    .COUT(_05603_),
    .SUM(_05604_));
 sky130_fd_sc_hd__ha_1 _11544_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[16] ),
    .COUT(_05605_),
    .SUM(_05606_));
 sky130_fd_sc_hd__ha_2 _11545_ (.A(\CPU_imm_a3[10] ),
    .B(_05541_),
    .COUT(_05607_),
    .SUM(_05608_));
 sky130_fd_sc_hd__ha_1 _11546_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[15] ),
    .COUT(_05609_),
    .SUM(_05610_));
 sky130_fd_sc_hd__ha_2 _11547_ (.A(\CPU_imm_a3[11] ),
    .B(_05546_),
    .COUT(_05611_),
    .SUM(_05612_));
 sky130_fd_sc_hd__ha_1 _11548_ (.A(\CPU_imm_a3[11] ),
    .B(\CPU_src1_value_a3[11] ),
    .COUT(_05613_),
    .SUM(_05614_));
 sky130_fd_sc_hd__ha_2 _11549_ (.A(\CPU_imm_a3[10] ),
    .B(_05551_),
    .COUT(_05615_),
    .SUM(_05616_));
 sky130_fd_sc_hd__ha_1 _11550_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[7] ),
    .COUT(_05617_),
    .SUM(_05618_));
 sky130_fd_sc_hd__ha_1 _11551_ (.A(\CPU_imm_a3[3] ),
    .B(_05556_),
    .COUT(_05619_),
    .SUM(_05620_));
 sky130_fd_sc_hd__ha_1 _11552_ (.A(\CPU_imm_a3[3] ),
    .B(\CPU_src1_value_a3[3] ),
    .COUT(_05621_),
    .SUM(_05622_));
 sky130_fd_sc_hd__ha_1 _11553_ (.A(\CPU_imm_a3[1] ),
    .B(_05511_),
    .COUT(_05623_),
    .SUM(_05624_));
 sky130_fd_sc_hd__ha_1 _11554_ (.A(\CPU_imm_a3[1] ),
    .B(\CPU_src1_value_a3[1] ),
    .COUT(_05625_),
    .SUM(_05626_));
 sky130_fd_sc_hd__ha_2 _11555_ (.A(_05627_),
    .B(\CPU_src1_value_a3[0] ),
    .COUT(_05628_),
    .SUM(_05629_));
 sky130_fd_sc_hd__ha_1 _11556_ (.A(\CPU_imm_a3[0] ),
    .B(\CPU_src1_value_a3[0] ),
    .COUT(_05630_),
    .SUM(_05631_));
 sky130_fd_sc_hd__ha_4 _11557_ (.A(\CPU_imm_a3[10] ),
    .B(_05523_),
    .COUT(_05632_),
    .SUM(_05633_));
 sky130_fd_sc_hd__ha_1 _11558_ (.A(\CPU_src1_value_a3[0] ),
    .B(_05634_),
    .COUT(_05635_),
    .SUM(_05636_));
 sky130_fd_sc_hd__ha_1 _11559_ (.A(\CPU_src1_value_a3[0] ),
    .B(\CPU_src2_value_a3[0] ),
    .COUT(_05637_),
    .SUM(_05638_));
 sky130_fd_sc_hd__ha_2 _11560_ (.A(\CPU_imm_a3[2] ),
    .B(_05639_),
    .COUT(_05640_),
    .SUM(_05641_));
 sky130_fd_sc_hd__ha_1 _11561_ (.A(\CPU_imm_a3[2] ),
    .B(\CPU_src1_value_a3[2] ),
    .COUT(_05642_),
    .SUM(_05643_));
 sky130_fd_sc_hd__ha_1 _11562_ (.A(_05639_),
    .B(\CPU_src2_value_a3[2] ),
    .COUT(_05644_),
    .SUM(_05645_));
 sky130_fd_sc_hd__ha_1 _11563_ (.A(\CPU_src1_value_a3[2] ),
    .B(\CPU_src2_value_a3[2] ),
    .COUT(_05646_),
    .SUM(_05647_));
 sky130_fd_sc_hd__ha_1 _11564_ (.A(\CPU_imm_a3[4] ),
    .B(_05648_),
    .COUT(_05649_),
    .SUM(_05650_));
 sky130_fd_sc_hd__ha_1 _11565_ (.A(\CPU_imm_a3[4] ),
    .B(\CPU_src1_value_a3[4] ),
    .COUT(_05651_),
    .SUM(_05652_));
 sky130_fd_sc_hd__ha_2 _11566_ (.A(_05648_),
    .B(\CPU_src2_value_a3[4] ),
    .COUT(_05653_),
    .SUM(_05654_));
 sky130_fd_sc_hd__ha_1 _11567_ (.A(\CPU_src1_value_a3[4] ),
    .B(\CPU_src2_value_a3[4] ),
    .COUT(_05655_),
    .SUM(_05656_));
 sky130_fd_sc_hd__ha_2 _11568_ (.A(\CPU_imm_a3[10] ),
    .B(_05657_),
    .COUT(_05658_),
    .SUM(_05659_));
 sky130_fd_sc_hd__ha_1 _11569_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[5] ),
    .COUT(_05660_),
    .SUM(_05661_));
 sky130_fd_sc_hd__ha_2 _11570_ (.A(_05657_),
    .B(\CPU_src2_value_a3[5] ),
    .COUT(_05662_),
    .SUM(_05663_));
 sky130_fd_sc_hd__ha_1 _11571_ (.A(\CPU_src1_value_a3[5] ),
    .B(\CPU_src2_value_a3[5] ),
    .COUT(_05664_),
    .SUM(_05665_));
 sky130_fd_sc_hd__ha_2 _11572_ (.A(\CPU_imm_a3[10] ),
    .B(_05666_),
    .COUT(_05667_),
    .SUM(_05668_));
 sky130_fd_sc_hd__ha_1 _11573_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[6] ),
    .COUT(_05669_),
    .SUM(_05670_));
 sky130_fd_sc_hd__ha_2 _11574_ (.A(_05666_),
    .B(\CPU_src2_value_a3[6] ),
    .COUT(_05671_),
    .SUM(_05672_));
 sky130_fd_sc_hd__ha_1 _11575_ (.A(\CPU_src1_value_a3[6] ),
    .B(\CPU_src2_value_a3[6] ),
    .COUT(_05673_),
    .SUM(_05674_));
 sky130_fd_sc_hd__ha_2 _11576_ (.A(\CPU_imm_a3[10] ),
    .B(_05675_),
    .COUT(_05676_),
    .SUM(_05677_));
 sky130_fd_sc_hd__ha_1 _11577_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[8] ),
    .COUT(_05678_),
    .SUM(_05679_));
 sky130_fd_sc_hd__ha_2 _11578_ (.A(_05675_),
    .B(\CPU_src2_value_a3[8] ),
    .COUT(_05680_),
    .SUM(_05681_));
 sky130_fd_sc_hd__ha_1 _11579_ (.A(\CPU_src1_value_a3[8] ),
    .B(\CPU_src2_value_a3[8] ),
    .COUT(_05682_),
    .SUM(_05683_));
 sky130_fd_sc_hd__ha_2 _11580_ (.A(\CPU_imm_a3[10] ),
    .B(_05684_),
    .COUT(_05685_),
    .SUM(_05686_));
 sky130_fd_sc_hd__ha_1 _11581_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[9] ),
    .COUT(_05687_),
    .SUM(_05688_));
 sky130_fd_sc_hd__ha_4 _11582_ (.A(_05684_),
    .B(\CPU_src2_value_a3[9] ),
    .COUT(_05689_),
    .SUM(_05690_));
 sky130_fd_sc_hd__ha_1 _11583_ (.A(\CPU_src1_value_a3[9] ),
    .B(\CPU_src2_value_a3[9] ),
    .COUT(_05691_),
    .SUM(_05692_));
 sky130_fd_sc_hd__ha_2 _11584_ (.A(\CPU_imm_a3[10] ),
    .B(_05693_),
    .COUT(_05694_),
    .SUM(_05695_));
 sky130_fd_sc_hd__ha_1 _11585_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[10] ),
    .COUT(_05696_),
    .SUM(_05697_));
 sky130_fd_sc_hd__ha_2 _11586_ (.A(_05693_),
    .B(\CPU_src2_value_a3[10] ),
    .COUT(_05698_),
    .SUM(_05699_));
 sky130_fd_sc_hd__ha_1 _11587_ (.A(\CPU_src1_value_a3[10] ),
    .B(\CPU_src2_value_a3[10] ),
    .COUT(_05700_),
    .SUM(_05701_));
 sky130_fd_sc_hd__ha_2 _11588_ (.A(\CPU_imm_a3[10] ),
    .B(_05702_),
    .COUT(_05703_),
    .SUM(_05704_));
 sky130_fd_sc_hd__ha_1 _11589_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[12] ),
    .COUT(_05705_),
    .SUM(_05706_));
 sky130_fd_sc_hd__ha_2 _11590_ (.A(_05702_),
    .B(\CPU_src2_value_a3[12] ),
    .COUT(_05707_),
    .SUM(_05708_));
 sky130_fd_sc_hd__ha_1 _11591_ (.A(\CPU_src1_value_a3[12] ),
    .B(\CPU_src2_value_a3[12] ),
    .COUT(_05709_),
    .SUM(_05710_));
 sky130_fd_sc_hd__ha_2 _11592_ (.A(\CPU_imm_a3[10] ),
    .B(_05711_),
    .COUT(_05712_),
    .SUM(_05713_));
 sky130_fd_sc_hd__ha_1 _11593_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[13] ),
    .COUT(_05714_),
    .SUM(_05715_));
 sky130_fd_sc_hd__ha_2 _11594_ (.A(_05711_),
    .B(\CPU_src2_value_a3[13] ),
    .COUT(_05716_),
    .SUM(_05717_));
 sky130_fd_sc_hd__ha_1 _11595_ (.A(\CPU_src1_value_a3[13] ),
    .B(\CPU_src2_value_a3[13] ),
    .COUT(_05718_),
    .SUM(_05719_));
 sky130_fd_sc_hd__ha_2 _11596_ (.A(\CPU_imm_a3[10] ),
    .B(_05720_),
    .COUT(_05721_),
    .SUM(_05722_));
 sky130_fd_sc_hd__ha_1 _11597_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[14] ),
    .COUT(_05723_),
    .SUM(_05724_));
 sky130_fd_sc_hd__ha_2 _11598_ (.A(_05720_),
    .B(\CPU_src2_value_a3[14] ),
    .COUT(_05725_),
    .SUM(_05726_));
 sky130_fd_sc_hd__ha_1 _11599_ (.A(\CPU_src1_value_a3[14] ),
    .B(\CPU_src2_value_a3[14] ),
    .COUT(_05727_),
    .SUM(_05728_));
 sky130_fd_sc_hd__ha_1 _11600_ (.A(_05602_),
    .B(\CPU_src2_value_a3[16] ),
    .COUT(_05729_),
    .SUM(_05730_));
 sky130_fd_sc_hd__ha_1 _11601_ (.A(\CPU_src1_value_a3[16] ),
    .B(\CPU_src2_value_a3[16] ),
    .COUT(_05731_),
    .SUM(_05732_));
 sky130_fd_sc_hd__ha_2 _11602_ (.A(_05597_),
    .B(\CPU_src2_value_a3[17] ),
    .COUT(_05733_),
    .SUM(_05734_));
 sky130_fd_sc_hd__ha_1 _11603_ (.A(\CPU_src1_value_a3[17] ),
    .B(\CPU_src2_value_a3[17] ),
    .COUT(_05735_),
    .SUM(_05736_));
 sky130_fd_sc_hd__ha_2 _11604_ (.A(\CPU_imm_a3[10] ),
    .B(_05737_),
    .COUT(_05738_),
    .SUM(_05739_));
 sky130_fd_sc_hd__ha_1 _11605_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[18] ),
    .COUT(_05740_),
    .SUM(_05741_));
 sky130_fd_sc_hd__ha_2 _11606_ (.A(_05737_),
    .B(\CPU_src2_value_a3[18] ),
    .COUT(_05742_),
    .SUM(_05743_));
 sky130_fd_sc_hd__ha_1 _11607_ (.A(\CPU_src1_value_a3[18] ),
    .B(\CPU_src2_value_a3[18] ),
    .COUT(_05744_),
    .SUM(_05745_));
 sky130_fd_sc_hd__ha_4 _11608_ (.A(\CPU_imm_a3[10] ),
    .B(_05746_),
    .COUT(_05747_),
    .SUM(_05748_));
 sky130_fd_sc_hd__ha_1 _11609_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[20] ),
    .COUT(_05749_),
    .SUM(_05750_));
 sky130_fd_sc_hd__ha_2 _11610_ (.A(_05746_),
    .B(\CPU_src2_value_a3[20] ),
    .COUT(_05751_),
    .SUM(_05752_));
 sky130_fd_sc_hd__ha_1 _11611_ (.A(\CPU_src1_value_a3[20] ),
    .B(\CPU_src2_value_a3[20] ),
    .COUT(_05753_),
    .SUM(_05754_));
 sky130_fd_sc_hd__ha_2 _11612_ (.A(\CPU_imm_a3[10] ),
    .B(_05755_),
    .COUT(_05756_),
    .SUM(_05757_));
 sky130_fd_sc_hd__ha_1 _11613_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[21] ),
    .COUT(_05758_),
    .SUM(_05759_));
 sky130_fd_sc_hd__ha_2 _11614_ (.A(_05755_),
    .B(\CPU_src2_value_a3[21] ),
    .COUT(_05760_),
    .SUM(_05761_));
 sky130_fd_sc_hd__ha_1 _11615_ (.A(\CPU_src1_value_a3[21] ),
    .B(\CPU_src2_value_a3[21] ),
    .COUT(_05762_),
    .SUM(_05763_));
 sky130_fd_sc_hd__ha_2 _11616_ (.A(\CPU_imm_a3[10] ),
    .B(_05764_),
    .COUT(_05765_),
    .SUM(_05766_));
 sky130_fd_sc_hd__ha_1 _11617_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[22] ),
    .COUT(_05767_),
    .SUM(_05768_));
 sky130_fd_sc_hd__ha_4 _11618_ (.A(_05764_),
    .B(\CPU_src2_value_a3[22] ),
    .COUT(_05769_),
    .SUM(_05770_));
 sky130_fd_sc_hd__ha_1 _11619_ (.A(\CPU_src1_value_a3[22] ),
    .B(\CPU_src2_value_a3[22] ),
    .COUT(_05771_),
    .SUM(_05772_));
 sky130_fd_sc_hd__ha_2 _11620_ (.A(_05584_),
    .B(\CPU_src2_value_a3[24] ),
    .COUT(_05773_),
    .SUM(_05774_));
 sky130_fd_sc_hd__ha_2 _11621_ (.A(\CPU_src1_value_a3[24] ),
    .B(\CPU_src2_value_a3[24] ),
    .COUT(_05775_),
    .SUM(_05776_));
 sky130_fd_sc_hd__ha_2 _11622_ (.A(_05579_),
    .B(\CPU_src2_value_a3[25] ),
    .COUT(_05777_),
    .SUM(_05778_));
 sky130_fd_sc_hd__ha_1 _11623_ (.A(\CPU_src1_value_a3[25] ),
    .B(\CPU_src2_value_a3[25] ),
    .COUT(_05779_),
    .SUM(_05780_));
 sky130_fd_sc_hd__ha_2 _11624_ (.A(\CPU_imm_a3[10] ),
    .B(_05781_),
    .COUT(_05782_),
    .SUM(_05783_));
 sky130_fd_sc_hd__ha_1 _11625_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[26] ),
    .COUT(_05784_),
    .SUM(_05785_));
 sky130_fd_sc_hd__ha_2 _11626_ (.A(_05781_),
    .B(\CPU_src2_value_a3[26] ),
    .COUT(_05786_),
    .SUM(_05787_));
 sky130_fd_sc_hd__ha_1 _11627_ (.A(\CPU_src1_value_a3[26] ),
    .B(\CPU_src2_value_a3[26] ),
    .COUT(_05788_),
    .SUM(_05789_));
 sky130_fd_sc_hd__ha_2 _11628_ (.A(_05570_),
    .B(\CPU_src2_value_a3[28] ),
    .COUT(_05790_),
    .SUM(_05791_));
 sky130_fd_sc_hd__ha_1 _11629_ (.A(\CPU_src1_value_a3[28] ),
    .B(\CPU_src2_value_a3[28] ),
    .COUT(_05792_),
    .SUM(_05793_));
 sky130_fd_sc_hd__ha_2 _11630_ (.A(_05565_),
    .B(\CPU_src2_value_a3[29] ),
    .COUT(_05794_),
    .SUM(_05795_));
 sky130_fd_sc_hd__ha_1 _11631_ (.A(\CPU_src1_value_a3[29] ),
    .B(\CPU_src2_value_a3[29] ),
    .COUT(_05796_),
    .SUM(_05797_));
 sky130_fd_sc_hd__ha_1 _11632_ (.A(\CPU_imm_a3[10] ),
    .B(_05798_),
    .COUT(_05799_),
    .SUM(_05800_));
 sky130_fd_sc_hd__ha_1 _11633_ (.A(\CPU_imm_a3[10] ),
    .B(\CPU_src1_value_a3[30] ),
    .COUT(_05801_),
    .SUM(_05802_));
 sky130_fd_sc_hd__ha_2 _11634_ (.A(_05798_),
    .B(\CPU_src2_value_a3[30] ),
    .COUT(_05803_),
    .SUM(_05804_));
 sky130_fd_sc_hd__ha_1 _11635_ (.A(\CPU_src1_value_a3[30] ),
    .B(\CPU_src2_value_a3[30] ),
    .COUT(_05805_),
    .SUM(_05806_));
 sky130_fd_sc_hd__ha_1 _11636_ (.A(\CPU_imm_a2[1] ),
    .B(\CPU_inc_pc_a2[1] ),
    .COUT(_05807_),
    .SUM(_05808_));
 sky130_fd_sc_hd__ha_1 _11637_ (.A(net161),
    .B(net1706),
    .COUT(_05809_),
    .SUM(_05810_));
 sky130_fd_sc_hd__ha_1 _11638_ (.A(net155),
    .B(net1730),
    .COUT(_05811_),
    .SUM(_05812_));
 sky130_fd_sc_hd__ha_1 _11639_ (.A(net152),
    .B(net1715),
    .COUT(_05813_),
    .SUM(_05814_));
 sky130_fd_sc_hd__ha_1 _11640_ (.A(net150),
    .B(net154),
    .COUT(_05815_),
    .SUM(\CPU_br_tgt_pc_a2[0] ));
 sky130_fd_sc_hd__ha_2 _11641_ (.A(\CPU_inc_pc_a1[2] ),
    .B(_05816_),
    .COUT(_05817_),
    .SUM(\CPU_inc_pc_a1[3] ));
 sky130_fd_sc_hd__ha_1 _11642_ (.A(\CPU_inc_pc_a1[2] ),
    .B(\CPU_imem_rd_addr_a1[1] ),
    .COUT(_05818_),
    .SUM(_05819_));
 sky130_fd_sc_hd__ha_4 _11643_ (.A(net1585),
    .B(_05816_),
    .COUT(_05820_),
    .SUM(_05821_));
 sky130_fd_sc_hd__ha_2 _11644_ (.A(\CPU_imem_rd_addr_a1[0] ),
    .B(\CPU_imem_rd_addr_a1[1] ),
    .COUT(_05822_),
    .SUM(_05823_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[0]$_DFF_P_  (.D(net144),
    .Q(net2),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[1]$_DFF_P_  (.D(net153),
    .Q(net3),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[2]$_DFF_P_  (.D(net158),
    .Q(net4),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[3]$_DFF_P_  (.D(net143),
    .Q(net5),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__dfxtp_2 \out[4]$_DFF_P_  (.D(net134),
    .Q(net6),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[5]$_DFF_P_  (.D(net140),
    .Q(net7),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[6]$_DFF_P_  (.D(net157),
    .Q(net8),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[7]$_DFF_P_  (.D(net137),
    .Q(net9),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[8]$_DFF_P_  (.D(net135),
    .Q(net10),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \out[9]$_DFF_P_  (.D(net142),
    .Q(net11),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2714 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(reset),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net2),
    .X(out[0]));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net3),
    .X(out[1]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(out[2]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .X(out[3]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .X(out[4]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .X(out[5]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .X(out[6]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(out[7]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(out[8]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(out[9]));
 sky130_fd_sc_hd__buf_8 wire12 (.A(_03684_),
    .X(net12));
 sky130_fd_sc_hd__buf_16 load_slew13 (.A(_03627_),
    .X(net13));
 sky130_fd_sc_hd__buf_8 load_slew14 (.A(_04742_),
    .X(net14));
 sky130_fd_sc_hd__buf_16 load_slew15 (.A(_04742_),
    .X(net15));
 sky130_fd_sc_hd__buf_8 load_slew16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_16 max_cap17 (.A(_04726_),
    .X(net17));
 sky130_fd_sc_hd__buf_8 wire18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_8 wire19 (.A(_04724_),
    .X(net19));
 sky130_fd_sc_hd__buf_6 load_slew20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_8 load_slew21 (.A(_04716_),
    .X(net21));
 sky130_fd_sc_hd__buf_16 load_slew22 (.A(_04716_),
    .X(net22));
 sky130_fd_sc_hd__buf_6 load_slew23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_8 wire24 (.A(_04713_),
    .X(net24));
 sky130_fd_sc_hd__buf_16 load_slew25 (.A(_04707_),
    .X(net25));
 sky130_fd_sc_hd__buf_8 wire26 (.A(_04707_),
    .X(net26));
 sky130_fd_sc_hd__buf_6 load_slew27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_8 load_slew28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_16 load_slew29 (.A(_04269_),
    .X(net29));
 sky130_fd_sc_hd__buf_16 max_cap30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_8 wire31 (.A(_04266_),
    .X(net31));
 sky130_fd_sc_hd__buf_8 load_slew32 (.A(_04264_),
    .X(net32));
 sky130_fd_sc_hd__buf_16 load_slew33 (.A(_04264_),
    .X(net33));
 sky130_fd_sc_hd__buf_8 load_slew34 (.A(_04245_),
    .X(net34));
 sky130_fd_sc_hd__buf_16 max_cap35 (.A(_04245_),
    .X(net35));
 sky130_fd_sc_hd__buf_8 load_slew36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_8 load_slew37 (.A(_04241_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 load_slew38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__buf_16 max_cap39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_16 load_slew40 (.A(_04234_),
    .X(net40));
 sky130_fd_sc_hd__buf_16 max_cap41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_8 wire42 (.A(_02404_),
    .X(net42));
 sky130_fd_sc_hd__buf_8 wire43 (.A(_02327_),
    .X(net43));
 sky130_fd_sc_hd__buf_8 wire44 (.A(_02327_),
    .X(net44));
 sky130_fd_sc_hd__buf_8 load_slew45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__buf_16 max_cap46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_6 wire47 (.A(_02324_),
    .X(net47));
 sky130_fd_sc_hd__buf_16 max_cap48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_16 max_cap49 (.A(_02252_),
    .X(net49));
 sky130_fd_sc_hd__buf_16 load_slew50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_16 max_cap51 (.A(_02169_),
    .X(net51));
 sky130_fd_sc_hd__buf_8 wire52 (.A(_02097_),
    .X(net52));
 sky130_fd_sc_hd__buf_8 load_slew53 (.A(_02097_),
    .X(net53));
 sky130_fd_sc_hd__buf_16 max_cap54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_8 wire55 (.A(_02018_),
    .X(net55));
 sky130_fd_sc_hd__buf_6 load_slew56 (.A(_02015_),
    .X(net56));
 sky130_fd_sc_hd__buf_6 load_slew57 (.A(_02015_),
    .X(net57));
 sky130_fd_sc_hd__buf_6 load_slew58 (.A(_02015_),
    .X(net58));
 sky130_fd_sc_hd__buf_6 wire59 (.A(net61),
    .X(net59));
 sky130_fd_sc_hd__buf_6 load_slew60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_6 load_slew61 (.A(_01939_),
    .X(net61));
 sky130_fd_sc_hd__buf_8 wire62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_16 max_cap63 (.A(_01934_),
    .X(net63));
 sky130_fd_sc_hd__buf_8 wire64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_16 max_cap65 (.A(_01861_),
    .X(net65));
 sky130_fd_sc_hd__buf_6 load_slew66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__buf_6 load_slew67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_6 load_slew68 (.A(_01858_),
    .X(net68));
 sky130_fd_sc_hd__buf_6 load_slew69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__buf_6 wire70 (.A(_01786_),
    .X(net70));
 sky130_fd_sc_hd__buf_8 load_slew71 (.A(_01786_),
    .X(net71));
 sky130_fd_sc_hd__buf_8 wire72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_16 load_slew73 (.A(_01782_),
    .X(net73));
 sky130_fd_sc_hd__buf_8 load_slew74 (.A(_01709_),
    .X(net74));
 sky130_fd_sc_hd__buf_8 load_slew75 (.A(_01709_),
    .X(net75));
 sky130_fd_sc_hd__buf_16 max_cap76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_16 load_slew77 (.A(_01628_),
    .X(net77));
 sky130_fd_sc_hd__buf_6 load_slew78 (.A(_01557_),
    .X(net78));
 sky130_fd_sc_hd__buf_8 wire79 (.A(_01557_),
    .X(net79));
 sky130_fd_sc_hd__buf_16 load_slew80 (.A(_01478_),
    .X(net80));
 sky130_fd_sc_hd__buf_16 max_cap81 (.A(_01478_),
    .X(net81));
 sky130_fd_sc_hd__buf_6 load_slew82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_6 wire83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_8 max_cap84 (.A(_01475_),
    .X(net84));
 sky130_fd_sc_hd__buf_8 load_slew85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_16 max_cap86 (.A(_01401_),
    .X(net86));
 sky130_fd_sc_hd__buf_16 max_cap87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_16 load_slew88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_8 load_slew89 (.A(_01319_),
    .X(net89));
 sky130_fd_sc_hd__buf_8 load_slew90 (.A(net92),
    .X(net90));
 sky130_fd_sc_hd__buf_6 load_slew91 (.A(_04700_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 max_cap92 (.A(_04700_),
    .X(net92));
 sky130_fd_sc_hd__buf_6 wire93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__buf_6 wire94 (.A(_04237_),
    .X(net94));
 sky130_fd_sc_hd__buf_8 load_slew95 (.A(_04237_),
    .X(net95));
 sky130_fd_sc_hd__buf_16 load_slew96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_16 load_slew97 (.A(_02586_),
    .X(net97));
 sky130_fd_sc_hd__buf_16 load_slew98 (.A(_02483_),
    .X(net98));
 sky130_fd_sc_hd__buf_8 max_cap99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_6 wire100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_8 max_cap101 (.A(_01177_),
    .X(net101));
 sky130_fd_sc_hd__buf_12 load_slew102 (.A(net107),
    .X(net102));
 sky130_fd_sc_hd__buf_16 load_slew103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_16 load_slew104 (.A(net107),
    .X(net104));
 sky130_fd_sc_hd__buf_16 load_slew105 (.A(net107),
    .X(net105));
 sky130_fd_sc_hd__buf_16 load_slew106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_16 load_slew107 (.A(CPU_reset_a4),
    .X(net107));
 sky130_fd_sc_hd__buf_16 load_slew108 (.A(CPU_reset_a3),
    .X(net108));
 sky130_fd_sc_hd__buf_16 load_slew109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_12 load_slew110 (.A(CPU_reset_a3),
    .X(net110));
 sky130_fd_sc_hd__conb_1 \CPU_is_bltu_a2$_DFF_P__111  (.LO(net111));
 sky130_fd_sc_hd__conb_1 \CPU_is_slt_a2$_DFF_P__112  (.LO(net112));
 sky130_fd_sc_hd__conb_1 \CPU_is_slti_a2$_DFF_P__113  (.LO(net113));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload9 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload10 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload11 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload12 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinv_4 clkload17 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__bufinv_16 clkload18 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__bufinv_16 clkload21 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__bufinv_16 clkload22 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload23 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload25 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__bufinv_16 clkload26 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_4 clkload27 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__bufinv_16 clkload28 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__inv_4 clkload29 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload30 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinv_2 clkload31 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__inv_6 clkload32 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload33 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload35 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload37 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload38 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload39 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload40 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload41 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload42 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload43 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload45 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload46 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload47 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkinv_2 clkload48 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_2 clkload49 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload50 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__bufinv_16 clkload51 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload52 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload53 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__bufinv_16 clkload55 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload56 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__inv_8 clkload57 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_4 clkload58 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__bufinv_16 clkload59 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload61 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload62 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload63 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload64 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload65 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__bufinv_16 clkload67 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload68 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__bufinv_16 clkload69 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload70 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload71 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkinv_2 clkload72 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload73 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload75 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload76 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload77 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload78 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload79 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload80 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload81 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload82 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload83 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload84 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload85 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload87 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload88 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__bufinv_16 clkload89 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload90 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload91 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload92 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload93 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_2 clkload94 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinv_4 clkload95 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__inv_4 clkload96 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload97 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__bufinv_16 clkload98 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload99 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_2 clkload100 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_1 clkload101 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload103 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload104 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload105 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload106 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload107 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload108 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload109 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload110 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_2 clkload111 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinv_2 clkload112 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload113 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload114 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\CPU_rd_a4[1] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(CPU_is_s_instr_a3),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(CPU_is_load_a2),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\CPU_rd_a2[1] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(CPU_is_addi_a2),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\CPU_rd_a2[3] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(CPU_reset_a2),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\CPU_rd_a2[0] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\CPU_rd_a4[3] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\CPU_inc_pc_a2[4] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\CPU_inc_pc_a2[5] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\CPU_rd_a4[2] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\CPU_rd_a4[4] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\CPU_rd_a4[0] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\CPU_inc_pc_a2[3] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\CPU_inc_pc_a2[2] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\CPU_rd_a2[2] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(CPU_is_s_instr_a2),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(CPU_rd_valid_a2),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(CPU_is_blt_a2),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\CPU_Xreg_value_a5[14][4] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\CPU_Xreg_value_a5[14][8] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\CPU_rd_a2[4] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\CPU_Xreg_value_a5[14][7] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\CPU_inc_pc_a1[0] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(CPU_is_add_a2),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\CPU_Xreg_value_a5[14][5] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(CPU_is_slt_a2),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\CPU_Xreg_value_a5[14][9] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\CPU_Xreg_value_a5[14][3] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\CPU_Xreg_value_a5[14][0] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\CPU_imm_a2[11] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(CPU_is_bltu_a2),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(CPU_valid_taken_br_a4),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\CPU_inc_pc_a1[1] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(CPU_is_slti_a2),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\CPU_imm_a2[0] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(CPU_dmem_rd_en_a4),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\CPU_imm_a2[4] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\CPU_Xreg_value_a5[14][1] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\CPU_inc_pc_a2[0] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\CPU_imm_a2[3] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\CPU_inc_pc_a2[1] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\CPU_Xreg_value_a5[14][6] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\CPU_Xreg_value_a5[14][2] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\CPU_imm_a2[1] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\CPU_src2_value_a3[3] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\CPU_imm_a2[2] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\CPU_src2_value_a3[24] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\CPU_src2_value_a3[26] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\CPU_src2_value_a3[1] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\CPU_Xreg_value_a4[14][6] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\CPU_Xreg_value_a4[14][4] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\CPU_src2_value_a3[30] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\CPU_Xreg_value_a4[14][2] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\CPU_src2_value_a3[2] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\CPU_src2_value_a3[4] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\CPU_Xreg_value_a4[14][1] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\CPU_Xreg_value_a4[14][9] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\CPU_src2_value_a3[25] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\CPU_rd_a3[4] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\CPU_src2_value_a3[29] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\CPU_src2_value_a3[10] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\CPU_rd_a3[0] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\CPU_src2_value_a3[14] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\CPU_imm_a2[10] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\CPU_Xreg_value_a4[14][5] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\CPU_src2_value_a3[12] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\CPU_imem_rd_addr_a1[1] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\CPU_src2_value_a3[22] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\CPU_src2_value_a3[0] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\CPU_src2_value_a3[17] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\CPU_Xreg_value_a4[14][3] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\CPU_src2_value_a3[9] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\CPU_src2_value_a3[5] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\CPU_src2_value_a3[7] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\CPU_src2_value_a3[11] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\CPU_Xreg_value_a4[14][0] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\CPU_imem_rd_addr_a1[0] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\CPU_src2_value_a3[27] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\CPU_src2_value_a3[19] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\CPU_Xreg_value_a4[14][8] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\CPU_src2_value_a3[28] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\CPU_src2_value_a3[6] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\CPU_src2_value_a3[16] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\CPU_src2_value_a3[20] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\CPU_src2_value_a3[21] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\CPU_src2_value_a3[18] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\CPU_Dmem_value_a5[4][24] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_00336_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\CPU_Dmem_value_a5[9][20] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_00492_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\CPU_Dmem_value_a5[5][20] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00364_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\CPU_Dmem_value_a5[6][21] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_00397_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\CPU_Dmem_value_a5[9][30] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_00503_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\CPU_Dmem_value_a5[14][4] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00186_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\CPU_src2_value_a3[23] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\CPU_Dmem_value_a5[7][27] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_00435_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\CPU_Dmem_value_a5[15][28] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00212_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\CPU_Dmem_value_a5[9][14] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_00485_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\CPU_Dmem_value_a5[6][14] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_00389_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\CPU_Dmem_value_a5[1][13] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_00228_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\CPU_Dmem_value_a5[6][11] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_00386_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\CPU_Dmem_value_a5[14][22] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00174_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\CPU_Dmem_value_a5[10][14] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_00037_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\CPU_Dmem_value_a5[3][24] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_00304_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\CPU_Dmem_value_a5[8][1] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_00459_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\CPU_Dmem_value_a5[6][4] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00410_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\CPU_Dmem_value_a5[3][20] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00300_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\CPU_Dmem_value_a5[9][12] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_00483_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\CPU_Dmem_value_a5[10][12] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00035_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\CPU_Dmem_value_a5[3][29] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_00309_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\CPU_Dmem_value_a5[9][16] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_00487_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\CPU_Dmem_value_a5[7][8] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_00446_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\CPU_Dmem_value_a5[13][14] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_00133_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\CPU_Dmem_value_a5[9][1] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_00491_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\CPU_Dmem_value_a5[12][25] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_00113_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\CPU_Dmem_value_a5[8][14] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_00453_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\CPU_Dmem_value_a5[14][26] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_00178_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\CPU_Dmem_value_a5[8][29] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_00469_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\CPU_Dmem_value_a5[1][14] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_00229_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\CPU_Dmem_value_a5[4][30] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_00343_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\CPU_Dmem_value_a5[8][25] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_00465_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\CPU_Dmem_value_a5[8][15] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_00454_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\CPU_Dmem_value_a5[6][12] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_00387_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\CPU_Dmem_value_a5[4][1] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_00331_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\CPU_Dmem_value_a5[3][10] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_00289_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\CPU_Dmem_value_a5[14][17] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_00168_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\CPU_Dmem_value_a5[3][21] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_00301_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\CPU_Dmem_value_a5[2][8] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_00286_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\CPU_Dmem_value_a5[4][26] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_00338_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\CPU_Dmem_value_a5[7][31] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_00440_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\CPU_Dmem_value_a5[6][24] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_00400_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\CPU_Dmem_value_a5[6][31] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_00408_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\CPU_Dmem_value_a5[3][26] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_00306_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\CPU_Dmem_value_a5[13][6] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00156_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\CPU_Dmem_value_a5[15][24] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_00208_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\CPU_Dmem_value_a5[7][13] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_00420_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\CPU_Dmem_value_a5[1][31] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_00248_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\CPU_Dmem_value_a5[0][11] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_00002_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\CPU_Dmem_value_a5[2][25] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_00273_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\CPU_Dmem_value_a5[2][20] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_00268_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\CPU_Dmem_value_a5[15][11] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_00194_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\CPU_Dmem_value_a5[7][20] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_00428_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\CPU_Dmem_value_a5[4][22] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_00334_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\CPU_Dmem_value_a5[15][14] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_00197_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\CPU_Dmem_value_a5[3][9] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_00319_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\CPU_Dmem_value_a5[0][14] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_00005_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\CPU_Dmem_value_a5[7][7] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_00445_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\CPU_Dmem_value_a5[14][7] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_00189_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\CPU_Dmem_value_a5[8][17] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_00456_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\CPU_Dmem_value_a5[7][11] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_00418_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\CPU_Dmem_value_a5[3][12] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_00291_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\CPU_Dmem_value_a5[3][4] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_00314_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\CPU_Dmem_value_a5[12][13] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_00100_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\CPU_Dmem_value_a5[6][18] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_00393_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\CPU_Dmem_value_a5[4][17] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_00328_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\CPU_Dmem_value_a5[11][20] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_00076_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\CPU_Dmem_value_a5[8][4] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_00474_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\CPU_Dmem_value_a5[6][10] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_00385_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\CPU_Dmem_value_a5[13][19] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_00138_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\CPU_Dmem_value_a5[10][18] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_00041_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\CPU_Dmem_value_a5[6][17] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_00392_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\CPU_Dmem_value_a5[11][13] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_00068_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\CPU_Dmem_value_a5[10][21] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_00045_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\CPU_Dmem_value_a5[14][10] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_00161_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\CPU_Dmem_value_a5[5][15] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_00358_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\CPU_Dmem_value_a5[11][12] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_00067_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\CPU_Dmem_value_a5[14][19] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_00170_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\CPU_Dmem_value_a5[6][25] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_00401_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\CPU_Dmem_value_a5[10][5] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_00059_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\CPU_Dmem_value_a5[5][24] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_00368_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\CPU_Dmem_value_a5[13][25] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_00145_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\CPU_Dmem_value_a5[2][17] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_00264_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\CPU_Dmem_value_a5[0][29] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_00021_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\CPU_Dmem_value_a5[0][12] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_00003_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\CPU_Dmem_value_a5[1][18] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_00233_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\CPU_Dmem_value_a5[15][19] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_00202_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\CPU_Dmem_value_a5[9][29] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_00501_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\CPU_Dmem_value_a5[7][9] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_00447_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\CPU_Dmem_value_a5[3][11] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_00290_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\CPU_Dmem_value_a5[0][24] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_00016_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\CPU_Dmem_value_a5[5][6] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_00380_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\CPU_Dmem_value_a5[0][1] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_00011_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\CPU_Dmem_value_a5[1][27] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_00243_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\CPU_Dmem_value_a5[1][16] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_00231_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\CPU_Dmem_value_a5[11][10] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_00065_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\CPU_Dmem_value_a5[2][16] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_00263_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\CPU_Dmem_value_a5[2][27] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_00275_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\CPU_Dmem_value_a5[0][2] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_00022_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\CPU_Dmem_value_a5[8][0] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_00448_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\CPU_Dmem_value_a5[8][21] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_00461_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\CPU_Dmem_value_a5[15][20] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_00204_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\CPU_Dmem_value_a5[11][30] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_00087_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\CPU_Dmem_value_a5[12][19] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_00106_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\CPU_Dmem_value_a5[11][19] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_00074_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\CPU_Dmem_value_a5[15][13] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_00196_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\CPU_Dmem_value_a5[6][28] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_00404_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\CPU_Dmem_value_a5[9][23] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_00495_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\CPU_Dmem_value_a5[9][4] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_00506_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\CPU_Dmem_value_a5[6][15] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_00390_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\CPU_Dmem_value_a5[4][16] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_00327_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\CPU_Dmem_value_a5[15][27] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_00211_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\CPU_Dmem_value_a5[14][5] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_00187_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\CPU_Dmem_value_a5[9][26] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_00498_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\CPU_Dmem_value_a5[13][26] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_00146_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\CPU_Dmem_value_a5[5][28] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_00372_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\CPU_Dmem_value_a5[8][11] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_00450_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\CPU_Dmem_value_a5[12][10] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_00097_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\CPU_src2_value_a3[8] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\CPU_Dmem_value_a5[7][25] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_00433_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\CPU_Dmem_value_a5[11][28] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_00084_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\CPU_Dmem_value_a5[3][28] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_00308_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\CPU_Dmem_value_a5[10][17] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_00040_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\CPU_Dmem_value_a5[8][19] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_00458_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\CPU_Dmem_value_a5[0][31] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_00024_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\CPU_Dmem_value_a5[12][27] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_00115_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\CPU_Dmem_value_a5[10][9] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_00063_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\CPU_Dmem_value_a5[10][10] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_00033_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\CPU_Dmem_value_a5[13][12] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_00131_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\CPU_Dmem_value_a5[12][17] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_00104_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\CPU_Dmem_value_a5[5][22] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_00366_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\CPU_Dmem_value_a5[5][13] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_00356_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\CPU_Dmem_value_a5[10][2] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_00054_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\CPU_Dmem_value_a5[2][24] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_00272_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\CPU_Dmem_value_a5[8][9] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_00479_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\CPU_Dmem_value_a5[0][15] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_00006_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\CPU_Dmem_value_a5[8][12] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_00451_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\CPU_Dmem_value_a5[12][21] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_00109_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\CPU_Dmem_value_a5[10][20] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_00044_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\CPU_Dmem_value_a5[10][25] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_00049_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\CPU_Dmem_value_a5[10][30] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_00055_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\CPU_Dmem_value_a5[2][4] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_00282_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\CPU_Dmem_value_a5[4][8] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_00350_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\CPU_Dmem_value_a5[0][5] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_00027_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\CPU_Dmem_value_a5[5][3] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_00377_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\CPU_Dmem_value_a5[10][8] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_00062_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\CPU_Dmem_value_a5[5][18] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_00361_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\CPU_Dmem_value_a5[4][29] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_00341_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\CPU_Dmem_value_a5[7][18] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_00425_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\CPU_Dmem_value_a5[0][10] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_00001_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\CPU_Dmem_value_a5[7][4] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_00442_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\CPU_Xreg_value_a4[14][7] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\CPU_Dmem_value_a5[13][1] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_00139_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\CPU_Dmem_value_a5[6][7] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_00413_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\CPU_Dmem_value_a5[15][4] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_00218_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\CPU_Dmem_value_a5[7][26] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_00434_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\CPU_Dmem_value_a5[2][3] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_00281_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\CPU_Dmem_value_a5[14][15] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_00166_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\CPU_Dmem_value_a5[12][4] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_00122_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\CPU_Dmem_value_a5[14][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_00160_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\CPU_Dmem_value_a5[7][29] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_00437_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\CPU_Dmem_value_a5[2][23] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_00271_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\CPU_Dmem_value_a5[1][8] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_00254_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\CPU_Dmem_value_a5[9][13] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_00484_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\CPU_Dmem_value_a5[11][17] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_00072_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\CPU_Dmem_value_a5[3][19] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_00298_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\CPU_Dmem_value_a5[10][11] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(_00034_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\CPU_Dmem_value_a5[9][7] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(_00509_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\CPU_Dmem_value_a5[0][13] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_00004_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\CPU_Dmem_value_a5[0][8] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(_00030_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\CPU_Dmem_value_a5[14][29] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_00181_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\CPU_Dmem_value_a5[0][19] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_00010_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\CPU_Dmem_value_a5[9][25] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_00497_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\CPU_Dmem_value_a5[3][3] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_00313_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\CPU_Dmem_value_a5[1][24] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_00240_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\CPU_Dmem_value_a5[12][0] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_00096_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\CPU_Dmem_value_a5[0][25] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_00017_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\CPU_Dmem_value_a5[10][24] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_00048_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\CPU_Dmem_value_a5[12][14] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_00101_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\CPU_Dmem_value_a5[11][29] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_00085_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\CPU_Dmem_value_a5[1][4] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_00250_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\CPU_Dmem_value_a5[9][19] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_00490_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\CPU_Dmem_value_a5[1][3] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_00249_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\CPU_Dmem_value_a5[9][18] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_00489_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\CPU_Dmem_value_a5[4][13] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_00324_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\CPU_Dmem_value_a5[1][17] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_00232_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\CPU_Dmem_value_a5[4][15] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_00326_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\CPU_Dmem_value_a5[14][21] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_00173_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\CPU_Dmem_value_a5[2][21] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_00269_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\CPU_Dmem_value_a5[4][23] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_00335_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\CPU_Dmem_value_a5[7][24] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_00432_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\CPU_Dmem_value_a5[7][15] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_00422_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\CPU_Dmem_value_a5[10][29] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_00053_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\CPU_Dmem_value_a5[8][7] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_00477_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\CPU_Dmem_value_a5[14][27] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_00179_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\CPU_Dmem_value_a5[7][5] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_00443_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\CPU_Dmem_value_a5[5][12] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_00355_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\CPU_Dmem_value_a5[8][18] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_00457_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\CPU_Dmem_value_a5[1][25] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_00241_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\CPU_src2_value_a3[15] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\CPU_Dmem_value_a5[2][26] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_00274_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\CPU_Dmem_value_a5[11][18] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_00073_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\CPU_Dmem_value_a5[5][17] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_00360_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\CPU_Dmem_value_a5[14][13] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_00164_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\CPU_Dmem_value_a5[4][14] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_00325_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\CPU_Dmem_value_a5[1][26] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_00242_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\CPU_Dmem_value_a5[1][10] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_00225_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\CPU_Dmem_value_a5[11][11] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_00066_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\CPU_Dmem_value_a5[7][22] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_00430_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\CPU_Dmem_value_a5[6][19] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_00394_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\CPU_Dmem_value_a5[11][31] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_00088_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\CPU_Dmem_value_a5[7][17] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_00424_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\CPU_Dmem_value_a5[12][20] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_00108_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\CPU_Dmem_value_a5[8][2] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_00470_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\CPU_Dmem_value_a5[12][7] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_00125_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\CPU_Dmem_value_a5[11][6] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_00092_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\CPU_Dmem_value_a5[11][15] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_00070_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\CPU_Dmem_value_a5[9][31] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_00504_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\CPU_Dmem_value_a5[7][21] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_00429_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\CPU_Dmem_value_a5[8][20] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_00460_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\CPU_Dmem_value_a5[9][24] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_00496_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\CPU_Dmem_value_a5[6][3] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_00409_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\CPU_Dmem_value_a5[1][30] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_00247_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\CPU_Dmem_value_a5[0][20] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_00012_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\CPU_Dmem_value_a5[7][28] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_00436_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\CPU_Dmem_value_a5[6][0] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_00384_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\CPU_Dmem_value_a5[5][7] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_00381_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\CPU_Dmem_value_a5[13][4] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_00154_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\CPU_Dmem_value_a5[13][17] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_00136_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\CPU_Dmem_value_a5[9][8] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_00510_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\CPU_Dmem_value_a5[15][26] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_00210_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\CPU_Dmem_value_a5[6][29] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_00405_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\CPU_Dmem_value_a5[14][23] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_00175_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\CPU_Dmem_value_a5[7][10] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_00417_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\CPU_Dmem_value_a5[6][26] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_00402_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\CPU_Dmem_value_a5[13][11] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_00130_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\CPU_Dmem_value_a5[11][8] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_00094_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\CPU_Dmem_value_a5[5][4] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_00378_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\CPU_Dmem_value_a5[3][13] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_00292_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\CPU_Dmem_value_a5[13][7] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_00157_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\CPU_Dmem_value_a5[11][21] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_00077_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\CPU_Dmem_value_a5[12][30] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_00119_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\CPU_Dmem_value_a5[6][20] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_00396_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\CPU_Dmem_value_a5[4][21] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_00333_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\CPU_Dmem_value_a5[5][11] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_00354_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\CPU_Dmem_value_a5[1][2] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_00246_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\CPU_Dmem_value_a5[2][14] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_00261_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\CPU_Dmem_value_a5[13][15] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_00134_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\CPU_Dmem_value_a5[14][18] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_00169_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\CPU_Dmem_value_a5[1][29] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_00245_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\CPU_Dmem_value_a5[12][18] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_00105_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\CPU_src2_value_a3[13] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\CPU_Dmem_value_a5[2][28] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_00276_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\CPU_Dmem_value_a5[14][6] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_00188_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\CPU_Dmem_value_a5[1][9] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(_00255_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\CPU_Dmem_value_a5[5][16] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(_00359_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\CPU_Dmem_value_a5[13][16] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_00135_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\CPU_Dmem_value_a5[14][28] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(_00180_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\CPU_Dmem_value_a5[2][0] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(_00256_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\CPU_Dmem_value_a5[7][16] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_00423_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\CPU_Dmem_value_a5[4][18] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_00329_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\CPU_Dmem_value_a5[15][7] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_00221_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\CPU_Dmem_value_a5[5][23] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_00367_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\CPU_Dmem_value_a5[15][8] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_00222_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\CPU_Dmem_value_a5[6][30] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_00407_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\CPU_Dmem_value_a5[0][4] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_00026_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\CPU_Dmem_value_a5[15][10] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_00193_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\CPU_Dmem_value_a5[1][15] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(_00230_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\CPU_Dmem_value_a5[2][18] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_00265_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\CPU_Dmem_value_a5[13][18] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_00137_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\CPU_Dmem_value_a5[8][13] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_00452_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\CPU_Dmem_value_a5[0][17] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_00008_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\CPU_Dmem_value_a5[8][22] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_00462_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\CPU_Dmem_value_a5[11][4] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_00090_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\CPU_Dmem_value_a5[6][22] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_00398_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\CPU_Dmem_value_a5[7][3] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_00441_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\CPU_inc_pc_a3[0] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_01029_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\CPU_Dmem_value_a5[0][28] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_00020_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\CPU_Dmem_value_a5[2][6] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_00284_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\CPU_Dmem_value_a5[1][12] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(_00227_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\CPU_Dmem_value_a5[4][7] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_00349_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\CPU_Dmem_value_a5[12][8] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_00126_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\CPU_Dmem_value_a5[8][8] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(_00478_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\CPU_Dmem_value_a5[5][21] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(_00365_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\CPU_Dmem_value_a5[2][11] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(_00258_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\CPU_Dmem_value_a5[5][30] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_00375_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\CPU_Dmem_value_a5[5][8] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_00382_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\CPU_Dmem_value_a5[2][30] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(_00279_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\CPU_Dmem_value_a5[0][23] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(_00015_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\CPU_Dmem_value_a5[14][12] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(_00163_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\CPU_Dmem_value_a5[12][29] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(_00117_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\CPU_Dmem_value_a5[14][24] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(_00176_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\CPU_Dmem_value_a5[14][11] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_00162_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\CPU_Dmem_value_a5[10][0] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(_00032_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\CPU_Dmem_value_a5[12][1] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(_00107_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\CPU_Dmem_value_a5[0][7] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(_00029_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\CPU_Dmem_value_a5[9][11] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_00482_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\CPU_Dmem_value_a5[2][12] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(_00259_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\CPU_Dmem_value_a5[9][28] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(_00500_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\CPU_Dmem_value_a5[5][25] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(_00369_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\CPU_Dmem_value_a5[1][21] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_00237_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\CPU_Dmem_value_a5[12][16] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_00103_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\CPU_Dmem_value_a5[15][9] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(_00223_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\CPU_Dmem_value_a5[11][2] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_00086_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\CPU_Dmem_value_a5[4][28] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_00340_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\CPU_Dmem_value_a5[13][22] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_00142_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\CPU_Dmem_value_a5[8][6] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(_00476_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\CPU_Dmem_value_a5[13][29] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(_00149_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\CPU_Dmem_value_a5[13][27] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_00147_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\CPU_Dmem_value_a5[2][15] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(_00262_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\CPU_Dmem_value_a5[10][23] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(_00047_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\CPU_Dmem_value_a5[4][4] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(_00346_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\CPU_Dmem_value_a5[12][28] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_00116_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\CPU_Dmem_value_a5[3][15] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_00294_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\CPU_imem_rd_addr_a1[2] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\CPU_Dmem_value_a5[15][12] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_00195_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\CPU_Dmem_value_a5[4][3] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_00345_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\CPU_Dmem_value_a5[9][5] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_00507_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\CPU_Dmem_value_a5[12][11] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00098_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\CPU_Dmem_value_a5[9][27] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_00499_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\CPU_Dmem_value_a5[0][21] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_00013_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\CPU_Dmem_value_a5[7][12] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_00419_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\CPU_Dmem_value_a5[6][8] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_00414_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\CPU_Dmem_value_a5[0][27] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_00019_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\CPU_Dmem_value_a5[6][16] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_00391_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\CPU_Dmem_value_a5[0][0] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_00000_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\CPU_Dmem_value_a5[10][27] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_00051_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\CPU_Dmem_value_a5[8][27] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_00467_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\CPU_Dmem_value_a5[2][7] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_00285_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\CPU_Dmem_value_a5[12][22] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_00110_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\CPU_Dmem_value_a5[15][30] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_00215_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\CPU_Dmem_value_a5[3][5] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_00315_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\CPU_Dmem_value_a5[6][27] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_00403_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\CPU_Dmem_value_a5[3][17] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_00296_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\CPU_Dmem_value_a5[11][14] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_00069_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\CPU_Dmem_value_a5[1][7] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_00253_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\CPU_Dmem_value_a5[3][8] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_00318_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\CPU_Dmem_value_a5[15][25] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_00209_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\CPU_Dmem_value_a5[15][22] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_00206_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\CPU_Dmem_value_a5[13][21] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_00141_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\CPU_Dmem_value_a5[4][11] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_00322_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\CPU_Dmem_value_a5[12][26] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_00114_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\CPU_Dmem_value_a5[1][1] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_00235_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\CPU_Dmem_value_a5[11][23] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_00079_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\CPU_Dmem_value_a5[8][28] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_00468_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\CPU_Dmem_value_a5[4][20] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_00332_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\CPU_Dmem_value_a5[0][6] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_00028_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\CPU_Dmem_value_a5[8][30] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_00471_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\CPU_Dmem_value_a5[3][18] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_00297_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\CPU_Dmem_value_a5[11][27] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_00083_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\CPU_Dmem_value_a5[9][6] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_00508_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\CPU_rd_a3[1] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\CPU_Dmem_value_a5[13][23] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(_00143_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\CPU_Dmem_value_a5[10][31] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_00056_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\CPU_Dmem_value_a5[3][23] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(_00303_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\CPU_Dmem_value_a5[6][6] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(_00412_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\CPU_Dmem_value_a5[10][13] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(_00036_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\CPU_Dmem_value_a5[4][19] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(_00330_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\CPU_Dmem_value_a5[13][31] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(_00152_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\CPU_Dmem_value_a5[5][26] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(_00370_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\CPU_src2_value_a3[31] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\CPU_Dmem_value_a5[8][23] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_00463_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\CPU_Dmem_value_a5[10][4] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_00058_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\CPU_Dmem_value_a5[12][23] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_00111_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\CPU_Dmem_value_a5[2][10] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_00257_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\CPU_Dmem_value_a5[1][11] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_00226_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\CPU_Dmem_value_a5[1][20] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_00236_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\CPU_Dmem_value_a5[9][22] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_00494_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\CPU_Dmem_value_a5[14][8] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_00190_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\CPU_Dmem_value_a5[5][1] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_00363_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\CPU_Dmem_value_a5[8][24] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_00464_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\CPU_Dmem_value_a5[1][28] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_00244_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\CPU_Dmem_value_a5[11][26] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_00082_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\CPU_Dmem_value_a5[10][16] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_00039_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\CPU_Dmem_value_a5[3][30] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_00311_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\CPU_Dmem_value_a5[10][26] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_00050_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\CPU_Dmem_value_a5[9][17] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_00488_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\CPU_Dmem_value_a5[10][6] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_00060_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\CPU_Dmem_value_a5[10][15] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_00038_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\CPU_Dmem_value_a5[15][5] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_00219_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\CPU_Dmem_value_a5[6][5] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_00411_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\CPU_Dmem_value_a5[1][5] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_00251_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\CPU_Dmem_value_a5[4][25] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_00337_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\CPU_Dmem_value_a5[2][29] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_00277_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\CPU_Dmem_value_a5[14][14] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_00165_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\CPU_Dmem_value_a5[4][10] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_00321_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\CPU_Dmem_value_a5[11][7] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_00093_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\CPU_Dmem_value_a5[15][29] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_00213_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\CPU_Dmem_value_a5[8][26] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_00466_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\CPU_Dmem_value_a5[2][22] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_00270_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\CPU_Dmem_value_a5[1][6] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_00252_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\CPU_Dmem_value_a5[11][16] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_00071_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\CPU_Dmem_value_a5[11][0] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_00064_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\CPU_Dmem_value_a5[15][21] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_00205_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\CPU_Dmem_value_a5[10][28] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_00052_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\CPU_Dmem_value_a5[2][13] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_00260_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\CPU_Dmem_value_a5[14][9] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_00191_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\CPU_Dmem_value_a5[8][10] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_00449_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\CPU_Dmem_value_a5[0][3] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_00025_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\CPU_Dmem_value_a5[13][5] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_00155_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\CPU_Dmem_value_a5[14][30] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_00183_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\CPU_Dmem_value_a5[3][16] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_00295_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\CPU_Dmem_value_a5[1][22] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_00238_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\CPU_Dmem_value_a5[5][29] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_00373_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\CPU_Dmem_value_a5[2][2] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_00278_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\CPU_Dmem_value_a5[5][31] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_00376_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\CPU_Dmem_value_a5[11][24] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_00080_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\CPU_Dmem_value_a5[2][19] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_00266_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\CPU_Dmem_value_a5[14][25] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_00177_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\CPU_Dmem_value_a5[13][28] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_00148_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\CPU_inc_pc_a3[3] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_01025_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\CPU_Dmem_value_a5[0][18] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_00009_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\CPU_Dmem_value_a5[3][25] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_00305_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\CPU_Dmem_value_a5[11][22] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_00078_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\CPU_Dmem_value_a5[15][23] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_00207_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\CPU_Dmem_value_a5[2][31] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_00280_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\CPU_Dmem_value_a5[15][15] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_00198_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\CPU_inc_pc_a3[1] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_01030_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\CPU_Dmem_value_a5[6][2] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_00406_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\CPU_Dmem_value_a5[10][7] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_00061_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\CPU_Dmem_value_a5[5][19] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_00362_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\CPU_Dmem_value_a5[3][14] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_00293_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\CPU_Dmem_value_a5[4][5] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_00347_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\CPU_Dmem_value_a5[9][21] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_00493_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\CPU_Dmem_value_a5[14][31] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_00184_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\CPU_Dmem_value_a5[13][30] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_00151_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\CPU_Dmem_value_a5[9][15] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_00486_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\CPU_Dmem_value_a5[4][0] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_00320_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\CPU_Xreg_value_a4[14][11] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\CPU_Dmem_value_a5[15][3] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(_00217_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\CPU_Dmem_value_a5[8][16] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(_00455_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\CPU_Dmem_value_a5[11][25] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(_00081_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\CPU_Dmem_value_a5[11][3] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(_00089_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\CPU_Dmem_value_a5[14][20] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_00172_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\CPU_Dmem_value_a5[3][22] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_00302_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\CPU_Dmem_value_a5[7][14] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(_00421_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\CPU_Dmem_value_a5[3][27] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(_00307_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\CPU_Dmem_value_a5[4][31] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(_00344_),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\CPU_Dmem_value_a5[4][2] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(_00342_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\CPU_Dmem_value_a5[10][1] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_00043_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\CPU_Dmem_value_a5[0][26] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(_00018_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\CPU_Dmem_value_a5[0][22] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(_00014_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\CPU_Dmem_value_a5[7][2] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(_00438_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\CPU_Dmem_value_a5[7][23] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(_00431_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\CPU_Dmem_value_a5[0][30] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(_00023_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\CPU_Dmem_value_a5[1][23] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(_00239_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\CPU_Dmem_value_a5[14][16] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(_00167_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\CPU_Xreg_value_a4[13][10] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\CPU_Dmem_value_a5[7][30] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_00439_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\CPU_Xreg_value_a4[11][13] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\CPU_Dmem_value_a5[13][24] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(_00144_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\CPU_Dmem_value_a5[6][13] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(_00388_),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\CPU_Dmem_value_a5[5][5] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(_00379_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\CPU_Dmem_value_a5[15][18] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(_00201_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\CPU_Dmem_value_a5[10][22] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(_00046_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\CPU_Xreg_value_a4[9][6] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\CPU_rd_a3[2] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\CPU_Dmem_value_a5[12][12] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(_00099_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\CPU_Dmem_value_a5[3][2] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(_00310_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\CPU_Dmem_value_a5[12][24] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(_00112_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\CPU_Dmem_value_a5[13][13] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(_00132_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\CPU_Xreg_value_a4[2][13] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\CPU_Dmem_value_a5[1][0] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_00224_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\CPU_Dmem_value_a5[3][31] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_00312_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\CPU_Xreg_value_a4[3][11] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\CPU_Dmem_value_a5[3][7] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(_00317_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\CPU_Dmem_value_a5[12][15] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(_00102_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\CPU_Dmem_value_a5[7][6] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(_00444_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\CPU_Dmem_value_a5[15][17] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(_00200_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\CPU_Dmem_value_a5[10][3] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(_00057_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\CPU_Dmem_value_a5[13][10] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(_00129_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\CPU_Xreg_value_a4[4][13] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\CPU_Dmem_value_a5[15][31] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_00216_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\CPU_Xreg_value_a4[11][11] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\CPU_Xreg_value_a4[1][13] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\CPU_Dmem_value_a5[15][1] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_00203_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\CPU_Xreg_value_a4[1][5] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\CPU_Dmem_value_a5[9][0] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(_00480_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\CPU_Dmem_value_a5[6][23] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(_00399_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\CPU_Dmem_value_a5[15][6] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(_00220_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\CPU_Dmem_value_a5[7][19] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(_00426_),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\CPU_Dmem_value_a5[13][20] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(_00140_),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\CPU_Xreg_value_a4[8][4] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(_00986_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\CPU_Xreg_value_a4[10][6] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\CPU_Dmem_value_a5[13][8] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_00158_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\CPU_Dmem_value_a5[2][9] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_00287_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\CPU_Dmem_value_a5[8][31] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_00472_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\CPU_Dmem_value_a5[4][6] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_00348_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\CPU_Dmem_value_a5[8][3] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_00473_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\CPU_Dmem_value_a5[0][16] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_00007_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\CPU_Dmem_value_a5[3][6] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_00316_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\CPU_Dmem_value_a5[8][5] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_00475_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\CPU_Xreg_value_a4[4][4] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_00858_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\CPU_Xreg_value_a4[3][24] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\CPU_Dmem_value_a5[7][1] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(_00427_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\CPU_Xreg_value_a4[2][11] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\CPU_Dmem_value_a5[11][5] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_00091_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\CPU_Xreg_value_a4[4][11] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\CPU_Xreg_value_a4[9][13] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\CPU_Dmem_value_a5[6][1] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_00395_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\CPU_Dmem_value_a5[5][14] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_00357_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\CPU_Xreg_value_a4[3][4] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_00826_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\CPU_Xreg_value_a4[8][13] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\CPU_Xreg_value_a4[8][10] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\CPU_Xreg_value_a4[3][13] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\CPU_Dmem_value_a5[1][19] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(_00234_),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\CPU_Xreg_value_a4[7][11] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\CPU_Xreg_value_a4[1][11] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\CPU_Dmem_value_a5[5][2] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(_00374_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\CPU_Dmem_value_a5[12][9] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(_00127_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\CPU_Dmem_value_a5[9][10] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(_00481_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\CPU_Xreg_value_a4[13][4] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(_00666_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\CPU_Dmem_value_a5[2][5] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(_00283_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\CPU_Xreg_value_a4[12][26] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\CPU_Dmem_value_a5[12][6] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_00124_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\CPU_Dmem_value_a5[15][0] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_00192_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\CPU_Dmem_value_a5[10][19] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_00042_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\CPU_Dmem_value_a5[11][1] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_00075_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\CPU_Dmem_value_a5[15][16] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_00199_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\CPU_Xreg_value_a4[4][26] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\CPU_Xreg_value_a4[6][6] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(CPU_reset_a1),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\CPU_Xreg_value_a4[2][24] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\CPU_Xreg_value_a4[12][24] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\CPU_Xreg_value_a4[11][4] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(_00602_),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\CPU_Dmem_value_a5[12][2] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(_00118_),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\CPU_Dmem_value_a5[14][2] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(_00182_),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\CPU_Xreg_value_a4[2][26] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\CPU_Xreg_value_a4[10][5] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\CPU_Xreg_value_a4[11][6] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\CPU_Xreg_value_a4[3][26] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\CPU_Xreg_value_a4[10][4] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(_00570_),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\CPU_Dmem_value_a5[5][9] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(_00383_),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\CPU_Dmem_value_a5[12][3] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(_00121_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\CPU_Xreg_value_a4[5][6] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\CPU_Xreg_value_a4[12][13] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\CPU_Xreg_value_a4[15][13] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\CPU_Xreg_value_a4[12][10] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\CPU_Dmem_value_a5[7][0] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(_00416_),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\CPU_Xreg_value_a4[5][4] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(_00890_),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\CPU_Xreg_value_a4[11][24] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\CPU_Xreg_value_a4[1][24] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\CPU_Xreg_value_a4[6][4] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(_00922_),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\CPU_Xreg_value_a4[13][6] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\CPU_Dmem_value_a5[13][9] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_00159_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\CPU_Xreg_value_a4[7][5] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\CPU_Dmem_value_a5[3][1] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(_00299_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\CPU_Dmem_value_a5[13][0] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(_00128_),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\CPU_Xreg_value_a4[7][10] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\CPU_Dmem_value_a5[4][27] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_00339_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\CPU_Xreg_value_a4[3][5] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\CPU_Dmem_value_a5[14][3] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(_00185_),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\CPU_Dmem_value_a5[2][1] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(_00267_),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\CPU_Dmem_value_a5[4][12] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(_00323_),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\CPU_rd_a3[3] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\CPU_Dmem_value_a5[13][3] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_00153_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\CPU_Xreg_value_a4[0][29] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\CPU_Xreg_value_a4[14][10] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\CPU_Xreg_value_a4[8][11] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\CPU_Xreg_value_a4[0][14] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\CPU_Xreg_value_a4[8][26] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\CPU_Xreg_value_a4[15][4] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(_00730_),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\CPU_Dmem_value_a5[5][27] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(_00371_),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\CPU_Xreg_value_a4[15][5] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\CPU_Xreg_value_a4[2][4] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_00794_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\CPU_Xreg_value_a4[15][10] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\CPU_Xreg_value_a4[0][25] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\CPU_Xreg_value_a4[1][4] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_00762_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\CPU_Xreg_value_a4[7][26] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\CPU_Xreg_value_a4[11][5] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\CPU_Xreg_value_a4[5][11] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\CPU_Xreg_value_a4[12][4] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(_00634_),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\CPU_Xreg_value_a4[1][10] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\CPU_Xreg_value_a4[7][6] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\CPU_Xreg_value_a4[1][6] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\CPU_Xreg_value_a4[4][24] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\CPU_imem_rd_addr_a1[3] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\CPU_Xreg_value_a4[0][10] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\CPU_Xreg_value_a4[5][5] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\CPU_Xreg_value_a4[15][6] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\CPU_Xreg_value_a4[4][6] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\CPU_Xreg_value_a4[12][6] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\CPU_Xreg_value_a4[2][10] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\CPU_Xreg_value_a4[7][13] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\CPU_Xreg_value_a4[5][10] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\CPU_Dmem_value_a5[14][1] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_00171_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\CPU_br_tgt_pc_a3[2] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_04192_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\CPU_Xreg_value_a4[2][5] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\CPU_Xreg_value_a4[2][6] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\CPU_Xreg_value_a4[11][10] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\CPU_Xreg_value_a4[0][15] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\CPU_Xreg_value_a4[3][10] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\CPU_Xreg_value_a4[14][24] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\CPU_Dmem_value_a5[5][10] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_00353_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\CPU_Xreg_value_a4[0][16] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\CPU_Dmem_value_a5[5][0] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(_00352_),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(\CPU_Xreg_value_a4[13][11] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\CPU_Dmem_value_a5[15][2] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_00214_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\CPU_Xreg_value_a4[6][5] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\CPU_Xreg_value_a4[7][24] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\CPU_Xreg_value_a4[10][11] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\CPU_Dmem_value_a5[9][3] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(_00505_),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\CPU_Xreg_value_a4[12][9] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\CPU_Xreg_value_a4[5][24] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\CPU_Xreg_value_a4[8][5] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\CPU_Xreg_value_a4[15][24] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\CPU_Xreg_value_a4[9][4] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(_01018_),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\CPU_Dmem_value_a5[11][9] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(_00095_),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\CPU_Xreg_value_a4[8][24] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\CPU_Xreg_value_a4[10][9] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\CPU_Xreg_value_a4[1][26] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\CPU_Xreg_value_a4[13][5] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\CPU_Xreg_value_a4[15][11] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\CPU_Xreg_value_a4[15][26] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\CPU_Xreg_value_a4[11][26] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\CPU_Xreg_value_a4[7][4] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_00954_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\CPU_Xreg_value_a4[12][11] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\CPU_Dmem_value_a5[9][2] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(_00502_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\CPU_Xreg_value_a4[8][6] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\CPU_Dmem_value_a5[12][5] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_00123_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\CPU_Xreg_value_a4[9][26] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\CPU_Xreg_value_a4[4][10] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\CPU_Dmem_value_a5[13][2] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_00150_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\CPU_Xreg_value_a4[9][8] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\CPU_Xreg_value_a4[6][15] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\CPU_Dmem_value_a5[9][9] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_00511_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\CPU_Xreg_value_a4[5][26] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\CPU_Xreg_value_a4[15][8] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\CPU_Xreg_value_a4[10][10] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\CPU_Xreg_value_a4[5][13] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\CPU_Xreg_value_a4[9][11] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\CPU_Xreg_value_a4[3][6] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\CPU_Xreg_value_a4[14][26] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\CPU_Xreg_value_a4[14][13] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\CPU_Dmem_value_a5[4][9] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_00351_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\CPU_Xreg_value_a4[6][8] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\CPU_Xreg_value_a4[9][14] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\CPU_Xreg_value_a4[9][10] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\CPU_Xreg_value_a4[12][15] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\CPU_Xreg_value_a4[12][7] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\CPU_Xreg_value_a4[4][15] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\CPU_Xreg_value_a4[7][9] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(\CPU_Xreg_value_a4[14][15] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\CPU_Xreg_value_a4[13][24] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\CPU_Xreg_value_a4[5][14] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\CPU_Xreg_value_a4[8][9] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\CPU_Xreg_value_a4[9][24] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\CPU_Xreg_value_a4[3][14] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\CPU_Xreg_value_a4[6][16] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\CPU_Xreg_value_a4[8][14] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\CPU_Xreg_value_a4[7][15] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\CPU_Xreg_value_a4[13][16] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\CPU_Dmem_value_a5[0][9] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(_00031_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\CPU_Xreg_value_a4[4][9] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\CPU_Xreg_value_a4[3][16] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\CPU_Xreg_value_a4[6][10] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\CPU_Xreg_value_a4[4][8] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(\CPU_Xreg_value_a4[3][7] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\CPU_Xreg_value_a4[9][5] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\CPU_Xreg_value_a4[6][11] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\CPU_Xreg_value_a4[9][16] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\CPU_Xreg_value_a4[13][13] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\CPU_Xreg_value_a4[3][9] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\CPU_Xreg_value_a4[7][7] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\CPU_Xreg_value_a4[11][14] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\CPU_Xreg_value_a4[9][15] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\CPU_Xreg_value_a4[1][9] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\CPU_Xreg_value_a4[2][14] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\CPU_Xreg_value_a4[14][16] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\CPU_Xreg_value_a4[15][15] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\CPU_Xreg_value_a4[3][8] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\CPU_Xreg_value_a4[15][16] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\CPU_Xreg_value_a4[10][14] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\CPU_Xreg_value_a4[12][16] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\CPU_Xreg_value_a4[10][13] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\CPU_Xreg_value_a4[10][24] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\CPU_Xreg_value_a4[7][8] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\CPU_Xreg_value_a4[6][24] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\CPU_Xreg_value_a4[5][0] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\CPU_Xreg_value_a4[0][19] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\CPU_Xreg_value_a4[4][2] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\CPU_Xreg_value_a4[13][26] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\CPU_Xreg_value_a4[15][9] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\CPU_Dmem_value_a5[3][0] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_00288_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\CPU_Xreg_value_a4[9][12] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\CPU_Xreg_value_a4[11][7] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\CPU_Xreg_value_a4[4][16] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\CPU_Xreg_value_a4[0][17] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\CPU_Xreg_value_a4[14][14] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\CPU_Xreg_value_a4[13][8] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\CPU_Xreg_value_a4[10][8] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\CPU_Dmem_value_a5[5][6] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\CPU_Xreg_value_a4[4][7] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\CPU_Xreg_value_a4[5][16] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\CPU_Xreg_value_a4[8][8] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\CPU_Xreg_value_a4[12][14] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\CPU_Xreg_value_a4[12][5] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\CPU_Xreg_value_a4[4][14] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\CPU_Xreg_value_a4[6][9] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\CPU_Xreg_value_a4[9][7] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\CPU_Xreg_value_a4[11][9] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\CPU_Xreg_value_a4[9][9] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\CPU_Xreg_value_a4[6][26] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\CPU_Xreg_value_a4[10][1] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\CPU_Xreg_value_a4[4][12] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\CPU_Xreg_value_a4[12][8] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\CPU_Xreg_value_a4[11][8] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\CPU_Xreg_value_a4[15][3] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\CPU_Xreg_value_a4[2][16] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\CPU_Xreg_value_a4[15][1] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\CPU_Xreg_value_a4[3][12] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\CPU_Xreg_value_a4[1][16] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\CPU_Xreg_value_a4[13][9] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\CPU_Xreg_value_a4[10][15] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\CPU_Xreg_value_a4[7][14] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\CPU_Xreg_value_a4[5][7] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\CPU_Xreg_value_a4[10][16] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\CPU_Xreg_value_a4[5][8] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\CPU_Xreg_value_a4[6][2] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\CPU_Xreg_value_a4[5][2] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\CPU_Xreg_value_a4[4][5] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\CPU_Xreg_value_a4[8][16] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\CPU_dmem_rd_data_a5[4] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\CPU_Xreg_value_a4[11][16] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\CPU_Xreg_value_a4[0][28] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\CPU_Xreg_value_a4[5][9] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\CPU_Xreg_value_a4[6][13] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\CPU_Xreg_value_a4[6][14] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\CPU_Xreg_value_a4[7][2] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\CPU_Xreg_value_a4[10][3] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\CPU_Xreg_value_a4[12][2] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\CPU_Xreg_value_a4[2][8] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\CPU_Xreg_value_a4[7][0] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\CPU_Xreg_value_a4[8][7] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\CPU_Xreg_value_a4[12][3] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\CPU_Xreg_value_a4[2][9] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\CPU_Xreg_value_a4[1][14] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\CPU_Xreg_value_a4[15][7] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\CPU_Xreg_value_a4[11][12] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\CPU_Xreg_value_a4[8][15] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\CPU_Xreg_value_a4[1][22] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\CPU_Xreg_value_a4[1][7] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\CPU_Xreg_value_a4[10][26] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\CPU_Xreg_value_a4[9][3] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\CPU_Xreg_value_a4[15][0] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\CPU_Xreg_value_a4[13][14] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\CPU_Xreg_value_a4[2][1] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\CPU_Xreg_value_a4[6][7] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(\CPU_Xreg_value_a4[2][7] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\CPU_Xreg_value_a4[8][21] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\CPU_Xreg_value_a4[12][12] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\CPU_Xreg_value_a4[15][14] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\CPU_Xreg_value_a4[3][0] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\CPU_Xreg_value_a4[11][27] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\CPU_Xreg_value_a4[1][0] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\CPU_Xreg_value_a4[8][3] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\CPU_Xreg_value_a4[6][12] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\CPU_Xreg_value_a4[11][1] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\CPU_Xreg_value_a4[7][21] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\CPU_Xreg_value_a4[3][1] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\CPU_Xreg_value_a4[12][1] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\CPU_Xreg_value_a4[13][2] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\CPU_Xreg_value_a4[13][7] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\CPU_Xreg_value_a4[1][12] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\CPU_Xreg_value_a4[8][27] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\CPU_Xreg_value_a4[13][15] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\CPU_Xreg_value_a4[1][8] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\CPU_Xreg_value_a4[15][17] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_00712_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\CPU_Xreg_value_a4[4][21] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\CPU_Xreg_value_a4[8][12] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\CPU_Xreg_value_a4[7][16] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\CPU_Xreg_value_a4[0][13] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\CPU_Xreg_value_a4[0][11] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\CPU_Xreg_value_a4[10][20] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(_00556_),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\CPU_Xreg_value_a4[11][3] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\CPU_Xreg_value_a4[7][29] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_00949_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\CPU_Xreg_value_a4[7][23] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\CPU_Xreg_value_a4[0][23] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\CPU_Xreg_value_a4[14][17] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_00680_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\CPU_Xreg_value_a4[9][0] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\CPU_Xreg_value_a4[10][27] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\CPU_Xreg_value_a4[6][23] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\CPU_Xreg_value_a4[3][3] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\CPU_Xreg_value_a4[4][27] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\CPU_Xreg_value_a4[10][23] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\CPU_Xreg_value_a4[0][3] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\CPU_Xreg_value_a4[8][1] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\CPU_Xreg_value_a4[15][27] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\CPU_Xreg_value_a4[5][12] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\CPU_Xreg_value_a4[5][20] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_00876_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\CPU_Xreg_value_a4[4][17] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_00840_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\CPU_Xreg_value_a4[9][29] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_01013_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\CPU_Xreg_value_a4[7][3] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\CPU_Xreg_value_a4[11][17] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(_00584_),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\CPU_Dmem_value_a5[12][31] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(_00120_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\CPU_Xreg_value_a4[13][29] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_00661_),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\CPU_Xreg_value_a4[7][1] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\CPU_Xreg_value_a4[8][20] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\CPU_Xreg_value_a4[2][21] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\CPU_Xreg_value_a4[7][20] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\CPU_Xreg_value_a4[15][23] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\CPU_Xreg_value_a4[0][24] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(\CPU_Xreg_value_a4[9][17] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(_01000_),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\CPU_Xreg_value_a4[5][21] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\CPU_Xreg_value_a4[13][12] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\CPU_Xreg_value_a4[8][29] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(_00981_),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\CPU_Xreg_value_a4[3][17] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(_00808_),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\CPU_Xreg_value_a4[4][23] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\CPU_Xreg_value_a4[15][2] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(\CPU_Xreg_value_a4[12][20] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\CPU_Xreg_value_a4[6][20] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\CPU_Xreg_value_a4[2][23] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\CPU_inc_pc_a3[4] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_04196_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(_01026_),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\CPU_Xreg_value_a4[14][29] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(_00693_),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(\CPU_Xreg_value_a4[2][2] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\CPU_Xreg_value_a4[10][29] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_00565_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\CPU_Xreg_value_a4[15][12] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\CPU_Xreg_value_a4[7][27] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\CPU_Xreg_value_a4[12][17] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_00616_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\CPU_Xreg_value_a4[2][15] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\CPU_imem_rd_addr_a1[2] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\CPU_Xreg_value_a4[9][2] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\CPU_Xreg_value_a4[0][26] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\CPU_Xreg_value_a4[4][3] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\CPU_Xreg_value_a4[10][17] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(_00552_),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\CPU_Xreg_value_a4[2][20] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\CPU_Xreg_value_a4[13][3] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\CPU_Xreg_value_a4[7][17] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(_00936_),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\CPU_Xreg_value_a4[1][2] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\CPU_Xreg_value_a4[11][21] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\CPU_inc_pc_a3[5] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(_04198_),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(_01027_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\CPU_Xreg_value_a4[8][23] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\CPU_imem_rd_addr_a1[0] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\CPU_Xreg_value_a4[1][20] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_00748_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\CPU_Xreg_value_a4[6][29] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\CPU_Xreg_value_a4[11][23] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\CPU_Xreg_value_a4[6][1] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\CPU_Xreg_value_a4[14][20] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(_00684_),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\CPU_Xreg_value_a4[15][29] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(_00725_),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\CPU_Xreg_value_a4[8][17] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(_00968_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\CPU_Xreg_value_a4[14][27] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\CPU_Xreg_value_a4[12][21] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\CPU_Xreg_value_a4[1][3] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\CPU_Xreg_value_a4[9][23] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\CPU_Xreg_value_a4[13][27] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\CPU_Xreg_value_a4[13][17] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_00648_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\CPU_Xreg_value_a4[6][27] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\CPU_Xreg_value_a4[5][17] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(_00872_),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\CPU_Xreg_value_a4[0][22] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\CPU_Xreg_value_a4[13][0] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\CPU_Xreg_value_a4[9][1] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\CPU_Xreg_value_a4[0][18] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\CPU_Xreg_value_a4[2][29] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\CPU_Xreg_value_a4[13][21] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\CPU_Xreg_value_a4[10][7] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\CPU_Xreg_value_a4[11][29] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\CPU_Xreg_value_a4[10][12] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\CPU_Xreg_value_a4[9][21] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\CPU_Xreg_value_a4[5][23] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\CPU_Xreg_value_a4[0][5] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\CPU_Xreg_value_a4[5][29] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(_00885_),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\CPU_Xreg_value_a4[10][2] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\CPU_Xreg_value_a4[14][21] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\CPU_Xreg_value_a4[12][27] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\CPU_Xreg_value_a4[13][1] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\CPU_Xreg_value_a4[1][27] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\CPU_Xreg_value_a4[4][20] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\CPU_Xreg_value_a4[3][2] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\CPU_Xreg_value_a4[11][15] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\CPU_Xreg_value_a4[11][20] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\CPU_Dmem_value_a5[6][9] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(_00415_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\CPU_Xreg_value_a4[1][1] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\CPU_Xreg_value_a4[1][29] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_00757_),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\CPU_Xreg_value_a4[2][12] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\CPU_Xreg_value_a4[15][21] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\CPU_Xreg_value_a4[3][29] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(_00821_),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\CPU_Xreg_value_a4[3][27] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\CPU_Xreg_value_a4[1][23] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\CPU_Xreg_value_a4[2][17] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(_00776_),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\CPU_Xreg_value_a4[5][15] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\CPU_Xreg_value_a4[1][17] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_00744_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\CPU_Xreg_value_a4[5][3] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\CPU_Xreg_value_a4[13][20] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(_00652_),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\CPU_Xreg_value_a4[10][21] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\CPU_Xreg_value_a4[4][1] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\CPU_Xreg_value_a4[9][27] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\CPU_Xreg_value_a4[11][0] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\CPU_Xreg_value_a4[15][20] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(_00716_),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\CPU_Xreg_value_a4[12][23] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\CPU_Xreg_value_a4[9][20] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_01004_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\CPU_Xreg_value_a4[5][27] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\CPU_Xreg_value_a4[5][1] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\CPU_Xreg_value_a4[6][17] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_00904_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\CPU_Xreg_value_a4[11][2] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\CPU_Xreg_value_a4[8][2] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\CPU_Xreg_value_a4[13][23] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\CPU_Xreg_value_a4[14][23] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\CPU_Xreg_value_a4[0][2] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(\CPU_Xreg_value_a4[2][3] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\CPU_Xreg_value_a4[6][3] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\CPU_Xreg_value_a4[0][27] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\CPU_Xreg_value_a4[1][15] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\CPU_Xreg_value_a4[0][21] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\CPU_Xreg_value_a4[6][21] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\CPU_Xreg_value_a4[0][4] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\CPU_Xreg_value_a4[0][8] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\CPU_Xreg_value_a4[0][20] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\CPU_Xreg_value_a4[0][1] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\CPU_Xreg_value_a4[3][21] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\CPU_Xreg_value_a4[0][9] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\CPU_Xreg_value_a4[0][0] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\CPU_Xreg_value_a4[12][29] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\CPU_Xreg_value_a4[3][20] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\CPU_Xreg_value_a4[1][21] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\CPU_Xreg_value_a4[0][31] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\CPU_Xreg_value_a4[0][12] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\CPU_Xreg_value_a4[0][6] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\CPU_Xreg_value_a4[4][29] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\CPU_Xreg_value_a4[2][27] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\CPU_Xreg_value_a4[3][23] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\CPU_Xreg_value_a4[0][7] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\CPU_Xreg_value_a4[0][30] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\CPU_Xreg_value_a4[14][12] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\CPU_Xreg_value_a4[12][25] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\CPU_pc_a2[5] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\CPU_br_tgt_pc_a2[5] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\CPU_Xreg_value_a4[1][25] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\CPU_Xreg_value_a4[15][25] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\CPU_Dmem_value_a5[12][9] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_05504_),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\CPU_Xreg_value_a4[7][25] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\CPU_Dmem_value_a5[13][8] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\CPU_Xreg_value_a4[8][25] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\CPU_Xreg_value_a4[2][25] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(\CPU_Xreg_value_a4[3][25] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\CPU_Xreg_value_a4[14][25] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\CPU_Xreg_value_a4[5][25] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\CPU_pc_a2[2] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\CPU_Xreg_value_a4[3][15] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\CPU_Dmem_value_a5[9][24] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\w_CPU_dmem_rd_data_a4[24] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\CPU_Xreg_value_a4[12][18] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\CPU_Xreg_value_a4[9][25] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\CPU_Xreg_value_a4[4][25] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\CPU_Xreg_value_a4[7][12] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\CPU_Xreg_value_a4[11][25] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\CPU_pc_a2[4] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\CPU_br_tgt_pc_a2[4] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\CPU_Xreg_value_a4[8][10] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(_04319_),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\CPU_Xreg_value_a4[3][25] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(_04980_),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(\CPU_Xreg_value_a4[13][25] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\CPU_Xreg_value_a4[10][25] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\CPU_Xreg_value_a4[1][25] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(_04521_),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_04522_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\CPU_Xreg_value_a4[9][28] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\CPU_Xreg_value_a4[11][18] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\CPU_Xreg_value_a4[3][18] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\CPU_Xreg_value_a4[12][31] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\CPU_pc_a2[3] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\CPU_Xreg_value_a4[4][18] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\CPU_Dmem_value_a5[2][11] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(\CPU_Xreg_value_a4[8][28] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\CPU_Xreg_value_a4[5][31] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\CPU_Xreg_value_a4[8][19] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\CPU_Xreg_value_a4[7][18] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\CPU_Xreg_value_a4[13][16] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\CPU_Xreg_value_a4[5][19] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\CPU_Xreg_value_a4[9][30] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\CPU_Xreg_value_a4[9][22] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\CPU_Xreg_value_a4[13][19] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\CPU_Xreg_value_a4[11][19] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\CPU_Xreg_value_a4[12][19] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\CPU_Xreg_value_a4[12][14] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_04374_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\CPU_Xreg_value_a4[6][19] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\CPU_Xreg_value_a4[3][19] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\CPU_Xreg_value_a4[10][28] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\CPU_Xreg_value_a4[3][30] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\CPU_Xreg_value_a4[7][19] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\CPU_Xreg_value_a4[10][19] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\CPU_Xreg_value_a4[15][31] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\CPU_Dmem_value_a5[2][22] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(_05331_),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\w_CPU_dmem_rd_data_a4[22] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\CPU_Xreg_value_a4[13][22] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\CPU_Xreg_value_a4[4][22] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\CPU_Xreg_value_a4[13][30] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\CPU_Xreg_value_a4[14][18] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\CPU_Xreg_value_a4[9][14] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_04838_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(_04839_),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\CPU_Xreg_value_a4[3][22] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\CPU_Xreg_value_a4[4][28] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\CPU_Xreg_value_a4[7][31] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\CPU_Xreg_value_a4[6][0] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\CPU_Xreg_value_a4[15][18] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\CPU_Xreg_value_a4[5][28] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\CPU_Xreg_value_a4[4][19] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\CPU_Xreg_value_a4[2][18] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\CPU_Xreg_value_a4[5][22] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\CPU_Xreg_value_a4[5][18] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\CPU_Xreg_value_a4[15][19] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\CPU_Xreg_value_a4[8][30] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\CPU_Xreg_value_a4[3][28] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\CPU_Xreg_value_a4[8][18] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\CPU_Xreg_value_a4[4][31] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\CPU_Xreg_value_a4[8][22] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\CPU_Xreg_value_a4[12][22] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\CPU_Xreg_value_a4[8][31] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\CPU_Xreg_value_a4[6][28] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\CPU_Xreg_value_a4[13][28] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\CPU_Xreg_value_a4[11][22] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\CPU_Xreg_value_a4[15][28] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\CPU_Xreg_value_a4[14][31] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\CPU_Dmem_value_a5[4][18] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_05282_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(_05285_),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\w_CPU_dmem_rd_data_a4[18] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\CPU_Xreg_value_a4[6][30] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\CPU_Xreg_value_a4[9][19] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\CPU_Xreg_value_a4[6][25] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\CPU_Xreg_value_a4[7][30] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\CPU_Xreg_value_a4[14][17] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\CPU_Xreg_value_a4[1][18] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\CPU_Xreg_value_a4[2][19] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\CPU_Xreg_value_a4[3][16] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(_04404_),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_04405_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\CPU_Xreg_value_a4[15][22] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\CPU_Xreg_value_a4[4][30] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\CPU_Xreg_value_a4[6][31] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\CPU_Xreg_value_a4[3][31] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\CPU_Xreg_value_a4[11][30] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\CPU_Xreg_value_a4[9][31] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\CPU_Xreg_value_a4[12][30] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\CPU_Xreg_value_a4[12][0] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\CPU_Xreg_value_a4[11][31] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\CPU_Xreg_value_a4[1][31] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\CPU_Xreg_value_a4[5][30] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\CPU_Xreg_value_a4[14][19] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\CPU_Xreg_value_a4[7][28] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\CPU_Xreg_value_a4[2][22] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\CPU_Xreg_value_a4[10][31] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\CPU_Xreg_value_a4[11][28] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\CPU_Xreg_value_a4[1][30] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\CPU_Xreg_value_a4[2][30] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\CPU_Xreg_value_a4[10][22] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\CPU_Xreg_value_a4[10][30] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\CPU_Xreg_value_a4[10][0] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\CPU_Dmem_value_a5[3][29] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\w_CPU_dmem_rd_data_a4[29] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\CPU_Xreg_value_a4[14][22] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\CPU_Xreg_value_a4[14][28] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\CPU_Xreg_value_a4[2][31] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\CPU_Xreg_value_a4[2][0] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\CPU_Xreg_value_a4[14][30] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\CPU_Xreg_value_a4[7][22] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\CPU_Xreg_value_a4[1][28] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\CPU_Dmem_value_a5[9][17] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(CPU_is_load_a3),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\CPU_Xreg_value_a4[4][0] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\CPU_imem_rd_addr_a1[3] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\CPU_Xreg_value_a4[15][30] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\CPU_Xreg_value_a4[10][18] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\CPU_Xreg_value_a4[9][18] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\CPU_Xreg_value_a4[1][19] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\CPU_Xreg_value_a4[13][18] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\CPU_Xreg_value_a4[12][28] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\CPU_Xreg_value_a4[8][0] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\CPU_Xreg_value_a4[6][22] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\CPU_Xreg_value_a4[6][18] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\CPU_Xreg_value_a4[13][31] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\CPU_Xreg_value_a4[2][28] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\CPU_Xreg_value_a4[4][18] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(_04425_),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\CPU_imem_rd_addr_a1[3] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\CPU_Xreg_value_a4[0][27] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\CPU_Xreg_value_a4[0][4] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\CPU_Xreg_value_a4[0][8] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\CPU_imem_rd_addr_a1[2] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\CPU_Xreg_value_a4[0][26] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\CPU_Xreg_value_a4[0][30] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\CPU_Xreg_value_a4[0][1] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\CPU_Xreg_value_a4[0][1] ),
    .X(net1855));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(CPU_reset_a1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04674_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_05141_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\w_CPU_dmem_rd_data_a4[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\w_CPU_dmem_rd_data_a4[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_01035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04958_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\w_CPU_dmem_rd_data_a4[14] ));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_780 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_911 ();
endmodule
